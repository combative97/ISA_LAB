LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Dadda_tree is PORT
(
	partial_p17_0,partial_p17_1,partial_p17_2,partial_p17_3,partial_p17_4,partial_p17_5,partial_p17_6,partial_p17_7,partial_p17_8,partial_p17_9,partial_p17_10,partial_p17_11,partial_p17_12,partial_p17_13,partial_p17_14,partial_p17_15,partial_p17_16 : IN std_logic_vector(63 downto 0);
	P : OUT std_logic_vector(63 downto 0)
);
END ENTITY;

Architecture beh of Dadda_tree is

component HA is
 
port( A,B : IN std_logic; 
     S,C : OUT std_logic); 
end component;

component FA is 
	port(A,B,Cin:in std_logic; 
		S,Cout:out std_logic); 
end component;


signal partial_p13_0,partial_p13_1,partial_p13_2,partial_p13_3,partial_p13_4,partial_p13_5,partial_p13_6,partial_p13_7,partial_p13_8,partial_p13_9,partial_p13_10,partial_p13_11,partial_p13_12 : std_logic_vector(63 downto 0);
signal partial_p9_0,partial_p9_1,partial_p9_2,partial_p9_3,partial_p9_4,partial_p9_5,partial_p9_6,partial_p9_7,partial_p9_8 : std_logic_vector (63 downto 0);
signal partial_p6_0,partial_p6_1,partial_p6_2,partial_p6_3,partial_p6_4,partial_p6_5 : std_logic_vector (63 downto 0);
signal partial_p4_0,partial_p4_1,partial_p4_2,partial_p4_3 : std_logic_vector (63 downto 0);
signal partial_p3_0,partial_p3_1,partial_p3_2 : std_logic_vector (63 downto 0);
signal partial_p2_0,partial_p2_1 : std_logic_vector (63 downto 0);
signal extra_carry : std_logic;
signal product : unsigned(63 downto 0);

begin

--LEVEL 1

partial_p13_0(0) <= partial_p17_0(0);
partial_p13_1(0) <= partial_p17_1(0);
partial_p13_2(0) <= partial_p17_2(0);
partial_p13_3(0) <= partial_p17_3(0);
partial_p13_4(0) <= partial_p17_4(0);
partial_p13_5(0) <= partial_p17_5(0);
partial_p13_6(0) <= partial_p17_6(0);
partial_p13_7(0) <= partial_p17_7(0);
partial_p13_8(0) <= partial_p17_8(0);
partial_p13_9(0) <= partial_p17_9(0);
partial_p13_10(0) <= partial_p17_10(0);
partial_p13_11(0) <= partial_p17_11(0);
partial_p13_12(0) <= partial_p17_12(0);
partial_p13_0(1) <= partial_p17_0(1);
partial_p13_1(1) <= partial_p17_1(1);
partial_p13_2(1) <= partial_p17_2(1);
partial_p13_3(1) <= partial_p17_3(1);
partial_p13_4(1) <= partial_p17_4(1);
partial_p13_5(1) <= partial_p17_5(1);
partial_p13_6(1) <= partial_p17_6(1);
partial_p13_7(1) <= partial_p17_7(1);
partial_p13_8(1) <= partial_p17_8(1);
partial_p13_9(1) <= partial_p17_9(1);
partial_p13_10(1) <= partial_p17_10(1);
partial_p13_11(1) <= partial_p17_11(1);
partial_p13_12(1) <= partial_p17_12(1);
partial_p13_0(2) <= partial_p17_0(2);
partial_p13_1(2) <= partial_p17_1(2);
partial_p13_2(2) <= partial_p17_2(2);
partial_p13_3(2) <= partial_p17_3(2);
partial_p13_4(2) <= partial_p17_4(2);
partial_p13_5(2) <= partial_p17_5(2);
partial_p13_6(2) <= partial_p17_6(2);
partial_p13_7(2) <= partial_p17_7(2);
partial_p13_8(2) <= partial_p17_8(2);
partial_p13_9(2) <= partial_p17_9(2);
partial_p13_10(2) <= partial_p17_10(2);
partial_p13_11(2) <= partial_p17_11(2);
partial_p13_12(2) <= partial_p17_12(2);
partial_p13_0(3) <= partial_p17_0(3);
partial_p13_1(3) <= partial_p17_1(3);
partial_p13_2(3) <= partial_p17_2(3);
partial_p13_3(3) <= partial_p17_3(3);
partial_p13_4(3) <= partial_p17_4(3);
partial_p13_5(3) <= partial_p17_5(3);
partial_p13_6(3) <= partial_p17_6(3);
partial_p13_7(3) <= partial_p17_7(3);
partial_p13_8(3) <= partial_p17_8(3);
partial_p13_9(3) <= partial_p17_9(3);
partial_p13_10(3) <= partial_p17_10(3);
partial_p13_11(3) <= partial_p17_11(3);
partial_p13_12(3) <= partial_p17_12(3);
partial_p13_0(4) <= partial_p17_0(4);
partial_p13_1(4) <= partial_p17_1(4);
partial_p13_2(4) <= partial_p17_2(4);
partial_p13_3(4) <= partial_p17_3(4);
partial_p13_4(4) <= partial_p17_4(4);
partial_p13_5(4) <= partial_p17_5(4);
partial_p13_6(4) <= partial_p17_6(4);
partial_p13_7(4) <= partial_p17_7(4);
partial_p13_8(4) <= partial_p17_8(4);
partial_p13_9(4) <= partial_p17_9(4);
partial_p13_10(4) <= partial_p17_10(4);
partial_p13_11(4) <= partial_p17_11(4);
partial_p13_12(4) <= partial_p17_12(4);
partial_p13_0(5) <= partial_p17_0(5);
partial_p13_1(5) <= partial_p17_1(5);
partial_p13_2(5) <= partial_p17_2(5);
partial_p13_3(5) <= partial_p17_3(5);
partial_p13_4(5) <= partial_p17_4(5);
partial_p13_5(5) <= partial_p17_5(5);
partial_p13_6(5) <= partial_p17_6(5);
partial_p13_7(5) <= partial_p17_7(5);
partial_p13_8(5) <= partial_p17_8(5);
partial_p13_9(5) <= partial_p17_9(5);
partial_p13_10(5) <= partial_p17_10(5);
partial_p13_11(5) <= partial_p17_11(5);
partial_p13_12(5) <= partial_p17_12(5);
partial_p13_0(6) <= partial_p17_0(6);
partial_p13_1(6) <= partial_p17_1(6);
partial_p13_2(6) <= partial_p17_2(6);
partial_p13_3(6) <= partial_p17_3(6);
partial_p13_4(6) <= partial_p17_4(6);
partial_p13_5(6) <= partial_p17_5(6);
partial_p13_6(6) <= partial_p17_6(6);
partial_p13_7(6) <= partial_p17_7(6);
partial_p13_8(6) <= partial_p17_8(6);
partial_p13_9(6) <= partial_p17_9(6);
partial_p13_10(6) <= partial_p17_10(6);
partial_p13_11(6) <= partial_p17_11(6);
partial_p13_12(6) <= partial_p17_12(6);
partial_p13_0(7) <= partial_p17_0(7);
partial_p13_1(7) <= partial_p17_1(7);
partial_p13_2(7) <= partial_p17_2(7);
partial_p13_3(7) <= partial_p17_3(7);
partial_p13_4(7) <= partial_p17_4(7);
partial_p13_5(7) <= partial_p17_5(7);
partial_p13_6(7) <= partial_p17_6(7);
partial_p13_7(7) <= partial_p17_7(7);
partial_p13_8(7) <= partial_p17_8(7);
partial_p13_9(7) <= partial_p17_9(7);
partial_p13_10(7) <= partial_p17_10(7);
partial_p13_11(7) <= partial_p17_11(7);
partial_p13_12(7) <= partial_p17_12(7);
partial_p13_0(8) <= partial_p17_0(8);
partial_p13_1(8) <= partial_p17_1(8);
partial_p13_2(8) <= partial_p17_2(8);
partial_p13_3(8) <= partial_p17_3(8);
partial_p13_4(8) <= partial_p17_4(8);
partial_p13_5(8) <= partial_p17_5(8);
partial_p13_6(8) <= partial_p17_6(8);
partial_p13_7(8) <= partial_p17_7(8);
partial_p13_8(8) <= partial_p17_8(8);
partial_p13_9(8) <= partial_p17_9(8);
partial_p13_10(8) <= partial_p17_10(8);
partial_p13_11(8) <= partial_p17_11(8);
partial_p13_12(8) <= partial_p17_12(8);
partial_p13_0(9) <= partial_p17_0(9);
partial_p13_1(9) <= partial_p17_1(9);
partial_p13_2(9) <= partial_p17_2(9);
partial_p13_3(9) <= partial_p17_3(9);
partial_p13_4(9) <= partial_p17_4(9);
partial_p13_5(9) <= partial_p17_5(9);
partial_p13_6(9) <= partial_p17_6(9);
partial_p13_7(9) <= partial_p17_7(9);
partial_p13_8(9) <= partial_p17_8(9);
partial_p13_9(9) <= partial_p17_9(9);
partial_p13_10(9) <= partial_p17_10(9);
partial_p13_11(9) <= partial_p17_11(9);
partial_p13_12(9) <= partial_p17_12(9);
partial_p13_0(10) <= partial_p17_0(10);
partial_p13_1(10) <= partial_p17_1(10);
partial_p13_2(10) <= partial_p17_2(10);
partial_p13_3(10) <= partial_p17_3(10);
partial_p13_4(10) <= partial_p17_4(10);
partial_p13_5(10) <= partial_p17_5(10);
partial_p13_6(10) <= partial_p17_6(10);
partial_p13_7(10) <= partial_p17_7(10);
partial_p13_8(10) <= partial_p17_8(10);
partial_p13_9(10) <= partial_p17_9(10);
partial_p13_10(10) <= partial_p17_10(10);
partial_p13_11(10) <= partial_p17_11(10);
partial_p13_12(10) <= partial_p17_12(10);
partial_p13_0(11) <= partial_p17_0(11);
partial_p13_1(11) <= partial_p17_1(11);
partial_p13_2(11) <= partial_p17_2(11);
partial_p13_3(11) <= partial_p17_3(11);
partial_p13_4(11) <= partial_p17_4(11);
partial_p13_5(11) <= partial_p17_5(11);
partial_p13_6(11) <= partial_p17_6(11);
partial_p13_7(11) <= partial_p17_7(11);
partial_p13_8(11) <= partial_p17_8(11);
partial_p13_9(11) <= partial_p17_9(11);
partial_p13_10(11) <= partial_p17_10(11);
partial_p13_11(11) <= partial_p17_11(11);
partial_p13_12(11) <= partial_p17_12(11);
partial_p13_0(12) <= partial_p17_0(12);
partial_p13_1(12) <= partial_p17_1(12);
partial_p13_2(12) <= partial_p17_2(12);
partial_p13_3(12) <= partial_p17_3(12);
partial_p13_4(12) <= partial_p17_4(12);
partial_p13_5(12) <= partial_p17_5(12);
partial_p13_6(12) <= partial_p17_6(12);
partial_p13_7(12) <= partial_p17_7(12);
partial_p13_8(12) <= partial_p17_8(12);
partial_p13_9(12) <= partial_p17_9(12);
partial_p13_10(12) <= partial_p17_10(12);
partial_p13_11(12) <= partial_p17_11(12);
partial_p13_12(12) <= partial_p17_12(12);
partial_p13_0(13) <= partial_p17_0(13);
partial_p13_1(13) <= partial_p17_1(13);
partial_p13_2(13) <= partial_p17_2(13);
partial_p13_3(13) <= partial_p17_3(13);
partial_p13_4(13) <= partial_p17_4(13);
partial_p13_5(13) <= partial_p17_5(13);
partial_p13_6(13) <= partial_p17_6(13);
partial_p13_7(13) <= partial_p17_7(13);
partial_p13_8(13) <= partial_p17_8(13);
partial_p13_9(13) <= partial_p17_9(13);
partial_p13_10(13) <= partial_p17_10(13);
partial_p13_11(13) <= partial_p17_11(13);
partial_p13_12(13) <= partial_p17_12(13);
partial_p13_0(14) <= partial_p17_0(14);
partial_p13_1(14) <= partial_p17_1(14);
partial_p13_2(14) <= partial_p17_2(14);
partial_p13_3(14) <= partial_p17_3(14);
partial_p13_4(14) <= partial_p17_4(14);
partial_p13_5(14) <= partial_p17_5(14);
partial_p13_6(14) <= partial_p17_6(14);
partial_p13_7(14) <= partial_p17_7(14);
partial_p13_8(14) <= partial_p17_8(14);
partial_p13_9(14) <= partial_p17_9(14);
partial_p13_10(14) <= partial_p17_10(14);
partial_p13_11(14) <= partial_p17_11(14);
partial_p13_12(14) <= partial_p17_12(14);
partial_p13_0(15) <= partial_p17_0(15);
partial_p13_1(15) <= partial_p17_1(15);
partial_p13_2(15) <= partial_p17_2(15);
partial_p13_3(15) <= partial_p17_3(15);
partial_p13_4(15) <= partial_p17_4(15);
partial_p13_5(15) <= partial_p17_5(15);
partial_p13_6(15) <= partial_p17_6(15);
partial_p13_7(15) <= partial_p17_7(15);
partial_p13_8(15) <= partial_p17_8(15);
partial_p13_9(15) <= partial_p17_9(15);
partial_p13_10(15) <= partial_p17_10(15);
partial_p13_11(15) <= partial_p17_11(15);
partial_p13_12(15) <= partial_p17_12(15);
partial_p13_0(16) <= partial_p17_0(16);
partial_p13_1(16) <= partial_p17_1(16);
partial_p13_2(16) <= partial_p17_2(16);
partial_p13_3(16) <= partial_p17_3(16);
partial_p13_4(16) <= partial_p17_4(16);
partial_p13_5(16) <= partial_p17_5(16);
partial_p13_6(16) <= partial_p17_6(16);
partial_p13_7(16) <= partial_p17_7(16);
partial_p13_8(16) <= partial_p17_8(16);
partial_p13_9(16) <= partial_p17_9(16);
partial_p13_10(16) <= partial_p17_10(16);
partial_p13_11(16) <= partial_p17_11(16);
partial_p13_12(16) <= partial_p17_12(16);
partial_p13_0(17) <= partial_p17_0(17);
partial_p13_1(17) <= partial_p17_1(17);
partial_p13_2(17) <= partial_p17_2(17);
partial_p13_3(17) <= partial_p17_3(17);
partial_p13_4(17) <= partial_p17_4(17);
partial_p13_5(17) <= partial_p17_5(17);
partial_p13_6(17) <= partial_p17_6(17);
partial_p13_7(17) <= partial_p17_7(17);
partial_p13_8(17) <= partial_p17_8(17);
partial_p13_9(17) <= partial_p17_9(17);
partial_p13_10(17) <= partial_p17_10(17);
partial_p13_11(17) <= partial_p17_11(17);
partial_p13_12(17) <= partial_p17_12(17);
partial_p13_0(18) <= partial_p17_0(18);
partial_p13_1(18) <= partial_p17_1(18);
partial_p13_2(18) <= partial_p17_2(18);
partial_p13_3(18) <= partial_p17_3(18);
partial_p13_4(18) <= partial_p17_4(18);
partial_p13_5(18) <= partial_p17_5(18);
partial_p13_6(18) <= partial_p17_6(18);
partial_p13_7(18) <= partial_p17_7(18);
partial_p13_8(18) <= partial_p17_8(18);
partial_p13_9(18) <= partial_p17_9(18);
partial_p13_10(18) <= partial_p17_10(18);
partial_p13_11(18) <= partial_p17_11(18);
partial_p13_12(18) <= partial_p17_12(18);
partial_p13_0(19) <= partial_p17_0(19);
partial_p13_1(19) <= partial_p17_1(19);
partial_p13_2(19) <= partial_p17_2(19);
partial_p13_3(19) <= partial_p17_3(19);
partial_p13_4(19) <= partial_p17_4(19);
partial_p13_5(19) <= partial_p17_5(19);
partial_p13_6(19) <= partial_p17_6(19);
partial_p13_7(19) <= partial_p17_7(19);
partial_p13_8(19) <= partial_p17_8(19);
partial_p13_9(19) <= partial_p17_9(19);
partial_p13_10(19) <= partial_p17_10(19);
partial_p13_11(19) <= partial_p17_11(19);
partial_p13_12(19) <= partial_p17_12(19);
partial_p13_0(20) <= partial_p17_0(20);
partial_p13_1(20) <= partial_p17_1(20);
partial_p13_2(20) <= partial_p17_2(20);
partial_p13_3(20) <= partial_p17_3(20);
partial_p13_4(20) <= partial_p17_4(20);
partial_p13_5(20) <= partial_p17_5(20);
partial_p13_6(20) <= partial_p17_6(20);
partial_p13_7(20) <= partial_p17_7(20);
partial_p13_8(20) <= partial_p17_8(20);
partial_p13_9(20) <= partial_p17_9(20);
partial_p13_10(20) <= partial_p17_10(20);
partial_p13_11(20) <= partial_p17_11(20);
partial_p13_12(20) <= partial_p17_12(20);
partial_p13_0(21) <= partial_p17_0(21);
partial_p13_1(21) <= partial_p17_1(21);
partial_p13_2(21) <= partial_p17_2(21);
partial_p13_3(21) <= partial_p17_3(21);
partial_p13_4(21) <= partial_p17_4(21);
partial_p13_5(21) <= partial_p17_5(21);
partial_p13_6(21) <= partial_p17_6(21);
partial_p13_7(21) <= partial_p17_7(21);
partial_p13_8(21) <= partial_p17_8(21);
partial_p13_9(21) <= partial_p17_9(21);
partial_p13_10(21) <= partial_p17_10(21);
partial_p13_11(21) <= partial_p17_11(21);
partial_p13_12(21) <= partial_p17_12(21);
partial_p13_0(22) <= partial_p17_0(22);
partial_p13_1(22) <= partial_p17_1(22);
partial_p13_2(22) <= partial_p17_2(22);
partial_p13_3(22) <= partial_p17_3(22);
partial_p13_4(22) <= partial_p17_4(22);
partial_p13_5(22) <= partial_p17_5(22);
partial_p13_6(22) <= partial_p17_6(22);
partial_p13_7(22) <= partial_p17_7(22);
partial_p13_8(22) <= partial_p17_8(22);
partial_p13_9(22) <= partial_p17_9(22);
partial_p13_10(22) <= partial_p17_10(22);
partial_p13_11(22) <= partial_p17_11(22);
partial_p13_12(22) <= partial_p17_12(22);
partial_p13_0(23) <= partial_p17_0(23);
partial_p13_1(23) <= partial_p17_1(23);
partial_p13_2(23) <= partial_p17_2(23);
partial_p13_3(23) <= partial_p17_3(23);
partial_p13_4(23) <= partial_p17_4(23);
partial_p13_5(23) <= partial_p17_5(23);
partial_p13_6(23) <= partial_p17_6(23);
partial_p13_7(23) <= partial_p17_7(23);
partial_p13_8(23) <= partial_p17_8(23);
partial_p13_9(23) <= partial_p17_9(23);
partial_p13_10(23) <= partial_p17_10(23);
partial_p13_11(23) <= partial_p17_11(23);
partial_p13_12(23) <= partial_p17_12(23);
HA_0 : HA port map(A=>partial_p17_0(24), B=>partial_p17_1(24), S=>partial_p13_0(24), C=>partial_p13_0(25));
partial_p13_1(24) <= partial_p17_2(24);
partial_p13_2(24) <= partial_p17_3(24);
partial_p13_3(24) <= partial_p17_4(24);
partial_p13_4(24) <= partial_p17_5(24);
partial_p13_5(24) <= partial_p17_6(24);
partial_p13_6(24) <= partial_p17_7(24);
partial_p13_7(24) <= partial_p17_8(24);
partial_p13_8(24) <= partial_p17_9(24);
partial_p13_9(24) <= partial_p17_10(24);
partial_p13_10(24) <= partial_p17_11(24);
partial_p13_11(24) <= partial_p17_12(24);
partial_p13_12(24) <= partial_p17_13(24);
HA_1 : HA port map(A=>partial_p17_0(25), B=>partial_p17_1(25), S=>partial_p13_1(25), C=>partial_p13_0(26));
partial_p13_2(25) <= partial_p17_2(25);
partial_p13_3(25) <= partial_p17_3(25);
partial_p13_4(25) <= partial_p17_4(25);
partial_p13_5(25) <= partial_p17_5(25);
partial_p13_6(25) <= partial_p17_6(25);
partial_p13_7(25) <= partial_p17_7(25);
partial_p13_8(25) <= partial_p17_8(25);
partial_p13_9(25) <= partial_p17_9(25);
partial_p13_10(25) <= partial_p17_10(25);
partial_p13_11(25) <= partial_p17_11(25);
partial_p13_12(25) <= partial_p17_12(25);
FA_0 : FA port map(A=>partial_p17_0(26), B=>partial_p17_1(26), Cin => partial_p17_2(26), S=>partial_p13_1(26), Cout=>partial_p13_0(27));
HA_2 : HA port map(A=>partial_p17_3(26), B=>partial_p17_4(26), S=>partial_p13_2(26), C=>partial_p13_1(27));
partial_p13_3(26) <= partial_p17_5(26);
partial_p13_4(26) <= partial_p17_6(26);
partial_p13_5(26) <= partial_p17_7(26);
partial_p13_6(26) <= partial_p17_8(26);
partial_p13_7(26) <= partial_p17_9(26);
partial_p13_8(26) <= partial_p17_10(26);
partial_p13_9(26) <= partial_p17_11(26);
partial_p13_10(26) <= partial_p17_12(26);
partial_p13_11(26) <= partial_p17_13(26);
partial_p13_12(26) <= partial_p17_14(26);
FA_1 : FA port map(A=>partial_p17_0(27), B=>partial_p17_1(27), Cin => partial_p17_2(27), S=>partial_p13_2(27), Cout=>partial_p13_0(28));
HA_3 : HA port map(A=>partial_p17_3(27), B=>partial_p17_4(27), S=>partial_p13_3(27), C=>partial_p13_1(28));
partial_p13_4(27) <= partial_p17_5(27);
partial_p13_5(27) <= partial_p17_6(27);
partial_p13_6(27) <= partial_p17_7(27);
partial_p13_7(27) <= partial_p17_8(27);
partial_p13_8(27) <= partial_p17_9(27);
partial_p13_9(27) <= partial_p17_10(27);
partial_p13_10(27) <= partial_p17_11(27);
partial_p13_11(27) <= partial_p17_12(27);
partial_p13_12(27) <= partial_p17_13(27);
FA_2 : FA port map(A=>partial_p17_0(28), B=>partial_p17_1(28), Cin => partial_p17_2(28), S=>partial_p13_2(28), Cout=>partial_p13_0(29));
FA_3 : FA port map(A=>partial_p17_3(28), B=>partial_p17_4(28), Cin => partial_p17_5(28), S=>partial_p13_3(28), Cout=>partial_p13_1(29));
HA_4 : HA port map(A=>partial_p17_6(28), B=>partial_p17_7(28), S=>partial_p13_4(28), C=>partial_p13_2(29));
partial_p13_5(28) <= partial_p17_8(28);
partial_p13_6(28) <= partial_p17_9(28);
partial_p13_7(28) <= partial_p17_10(28);
partial_p13_8(28) <= partial_p17_11(28);
partial_p13_9(28) <= partial_p17_12(28);
partial_p13_10(28) <= partial_p17_13(28);
partial_p13_11(28) <= partial_p17_14(28);
partial_p13_12(28) <= partial_p17_15(28);
FA_4 : FA port map(A=>partial_p17_0(29), B=>partial_p17_1(29), Cin => partial_p17_2(29), S=>partial_p13_3(29), Cout=>partial_p13_0(30));
FA_5 : FA port map(A=>partial_p17_3(29), B=>partial_p17_4(29), Cin => partial_p17_5(29), S=>partial_p13_4(29), Cout=>partial_p13_1(30));
HA_5 : HA port map(A=>partial_p17_6(29), B=>partial_p17_7(29), S=>partial_p13_5(29), C=>partial_p13_2(30));
partial_p13_6(29) <= partial_p17_8(29);
partial_p13_7(29) <= partial_p17_9(29);
partial_p13_8(29) <= partial_p17_10(29);
partial_p13_9(29) <= partial_p17_11(29);
partial_p13_10(29) <= partial_p17_12(29);
partial_p13_11(29) <= partial_p17_13(29);
partial_p13_12(29) <= partial_p17_14(29);
FA_6 : FA port map(A=>partial_p17_0(30), B=>partial_p17_1(30), Cin => partial_p17_2(30), S=>partial_p13_3(30), Cout=>partial_p13_0(31));
FA_7 : FA port map(A=>partial_p17_3(30), B=>partial_p17_4(30), Cin => partial_p17_5(30), S=>partial_p13_4(30), Cout=>partial_p13_1(31));
FA_8 : FA port map(A=>partial_p17_6(30), B=>partial_p17_7(30), Cin => partial_p17_8(30), S=>partial_p13_5(30), Cout=>partial_p13_2(31));
HA_6 : HA port map(A=>partial_p17_9(30), B=>partial_p17_10(30), S=>partial_p13_6(30), C=>partial_p13_3(31));
partial_p13_7(30) <= partial_p17_11(30);
partial_p13_8(30) <= partial_p17_12(30);
partial_p13_9(30) <= partial_p17_13(30);
partial_p13_10(30) <= partial_p17_14(30);
partial_p13_11(30) <= partial_p17_15(30);
partial_p13_12(30) <= partial_p17_16(30);
FA_9 : FA port map(A=>partial_p17_0(31), B=>partial_p17_1(31), Cin => partial_p17_2(31), S=>partial_p13_4(31), Cout=>partial_p13_0(32));
FA_10 : FA port map(A=>partial_p17_3(31), B=>partial_p17_4(31), Cin => partial_p17_5(31), S=>partial_p13_5(31), Cout=>partial_p13_1(32));
FA_11 : FA port map(A=>partial_p17_6(31), B=>partial_p17_7(31), Cin => partial_p17_8(31), S=>partial_p13_6(31), Cout=>partial_p13_2(32));
HA_7 : HA port map(A=>partial_p17_9(31), B=>partial_p17_10(31), S=>partial_p13_7(31), C=>partial_p13_3(32));
partial_p13_8(31) <= partial_p17_11(31);
partial_p13_9(31) <= partial_p17_12(31);
partial_p13_10(31) <= partial_p17_13(31);
partial_p13_11(31) <= partial_p17_14(31);
partial_p13_12(31) <= partial_p17_15(31);
FA_12 : FA port map(A=>partial_p17_0(32), B=>partial_p17_1(32), Cin => partial_p17_2(32), S=>partial_p13_4(32), Cout=>partial_p13_0(33));
FA_13 : FA port map(A=>partial_p17_3(32), B=>partial_p17_4(32), Cin => partial_p17_5(32), S=>partial_p13_5(32), Cout=>partial_p13_1(33));
FA_14 : FA port map(A=>partial_p17_6(32), B=>partial_p17_7(32), Cin => partial_p17_8(32), S=>partial_p13_6(32), Cout=>partial_p13_2(33));
FA_15 : FA port map(A=>partial_p17_9(32), B=>partial_p17_10(32), Cin => partial_p17_11(32), S=>partial_p13_7(32), Cout=>partial_p13_3(33));
partial_p13_8(32) <= partial_p17_12(32);
partial_p13_9(32) <= partial_p17_13(32);
partial_p13_10(32) <= partial_p17_14(32);
partial_p13_11(32) <= partial_p17_15(32);
partial_p13_12(32) <= partial_p17_16(32);
FA_16 : FA port map(A=>partial_p17_0(33), B=>partial_p17_1(33), Cin => partial_p17_2(33), S=>partial_p13_4(33), Cout=>partial_p13_0(34));
FA_17 : FA port map(A=>partial_p17_3(33), B=>partial_p17_4(33), Cin => partial_p17_5(33), S=>partial_p13_5(33), Cout=>partial_p13_1(34));
FA_18 : FA port map(A=>partial_p17_6(33), B=>partial_p17_7(33), Cin => partial_p17_8(33), S=>partial_p13_6(33), Cout=>partial_p13_2(34));
FA_19 : FA port map(A=>partial_p17_9(33), B=>partial_p17_10(33), Cin => partial_p17_11(33), S=>partial_p13_7(33), Cout=>partial_p13_3(34));
partial_p13_8(33) <= partial_p17_12(33);
partial_p13_9(33) <= partial_p17_13(33);
partial_p13_10(33) <= partial_p17_14(33);
partial_p13_11(33) <= partial_p17_15(33);
partial_p13_12(33) <= partial_p17_16(33);
FA_20 : FA port map(A=>partial_p17_0(34), B=>partial_p17_1(34), Cin => partial_p17_2(34), S=>partial_p13_4(34), Cout=>partial_p13_0(35));
FA_21 : FA port map(A=>partial_p17_3(34), B=>partial_p17_4(34), Cin => partial_p17_5(34), S=>partial_p13_5(34), Cout=>partial_p13_1(35));
FA_22 : FA port map(A=>partial_p17_6(34), B=>partial_p17_7(34), Cin => partial_p17_8(34), S=>partial_p13_6(34), Cout=>partial_p13_2(35));
FA_23 : FA port map(A=>partial_p17_9(34), B=>partial_p17_10(34), Cin => partial_p17_11(34), S=>partial_p13_7(34), Cout=>partial_p13_3(35));
partial_p13_8(34) <= partial_p17_12(34);
partial_p13_9(34) <= partial_p17_13(34);
partial_p13_10(34) <= partial_p17_14(34);
partial_p13_11(34) <= partial_p17_15(34);
partial_p13_12(34) <= partial_p17_16(34);
FA_24 : FA port map(A=>partial_p17_0(35), B=>partial_p17_1(35), Cin => partial_p17_2(35), S=>partial_p13_4(35), Cout=>partial_p13_0(36));
FA_25 : FA port map(A=>partial_p17_3(35), B=>partial_p17_4(35), Cin => partial_p17_5(35), S=>partial_p13_5(35), Cout=>partial_p13_1(36));
FA_26 : FA port map(A=>partial_p17_6(35), B=>partial_p17_7(35), Cin => partial_p17_8(35), S=>partial_p13_6(35), Cout=>partial_p13_2(36));
FA_27 : FA port map(A=>partial_p17_9(35), B=>partial_p17_10(35), Cin => partial_p17_11(35), S=>partial_p13_7(35), Cout=>partial_p13_3(36));
partial_p13_8(35) <= partial_p17_12(35);
partial_p13_9(35) <= partial_p17_13(35);
partial_p13_10(35) <= partial_p17_14(35);
partial_p13_11(35) <= partial_p17_15(35);
partial_p13_12(35) <= partial_p17_16(35);
FA_28 : FA port map(A=>partial_p17_0(36), B=>partial_p17_1(36), Cin => partial_p17_2(36), S=>partial_p13_4(36), Cout=>partial_p13_0(37));
FA_29 : FA port map(A=>partial_p17_3(36), B=>partial_p17_4(36), Cin => partial_p17_5(36), S=>partial_p13_5(36), Cout=>partial_p13_1(37));
FA_30 : FA port map(A=>partial_p17_6(36), B=>partial_p17_7(36), Cin => partial_p17_8(36), S=>partial_p13_6(36), Cout=>partial_p13_2(37));
HA_8 : HA port map(A=>partial_p17_9(36), B=>partial_p17_10(36), S=>partial_p13_7(36), C=>partial_p13_3(37));
partial_p13_8(36) <= partial_p17_11(36);
partial_p13_9(36) <= partial_p17_12(36);
partial_p13_10(36) <= partial_p17_13(36);
partial_p13_11(36) <= partial_p17_14(36);
partial_p13_12(36) <= partial_p17_15(36);
FA_31 : FA port map(A=>partial_p17_0(37), B=>partial_p17_1(37), Cin => partial_p17_2(37), S=>partial_p13_4(37), Cout=>partial_p13_0(38));
FA_32 : FA port map(A=>partial_p17_3(37), B=>partial_p17_4(37), Cin => partial_p17_5(37), S=>partial_p13_5(37), Cout=>partial_p13_1(38));
FA_33 : FA port map(A=>partial_p17_6(37), B=>partial_p17_7(37), Cin => partial_p17_8(37), S=>partial_p13_6(37), Cout=>partial_p13_2(38));
partial_p13_7(37) <= partial_p17_9(37);
partial_p13_8(37) <= partial_p17_10(37);
partial_p13_9(37) <= partial_p17_11(37);
partial_p13_10(37) <= partial_p17_12(37);
partial_p13_11(37) <= partial_p17_13(37);
partial_p13_12(37) <= partial_p17_14(37);
FA_34 : FA port map(A=>partial_p17_0(38), B=>partial_p17_1(38), Cin => partial_p17_2(38), S=>partial_p13_3(38), Cout=>partial_p13_0(39));
FA_35 : FA port map(A=>partial_p17_3(38), B=>partial_p17_4(38), Cin => partial_p17_5(38), S=>partial_p13_4(38), Cout=>partial_p13_1(39));
HA_9 : HA port map(A=>partial_p17_6(38), B=>partial_p17_7(38), S=>partial_p13_5(38), C=>partial_p13_2(39));
partial_p13_6(38) <= partial_p17_8(38);
partial_p13_7(38) <= partial_p17_9(38);
partial_p13_8(38) <= partial_p17_10(38);
partial_p13_9(38) <= partial_p17_11(38);
partial_p13_10(38) <= partial_p17_12(38);
partial_p13_11(38) <= partial_p17_13(38);
partial_p13_12(38) <= partial_p17_14(38);
FA_36 : FA port map(A=>partial_p17_0(39), B=>partial_p17_1(39), Cin => partial_p17_2(39), S=>partial_p13_3(39), Cout=>partial_p13_0(40));
FA_37 : FA port map(A=>partial_p17_3(39), B=>partial_p17_4(39), Cin => partial_p17_5(39), S=>partial_p13_4(39), Cout=>partial_p13_1(40));
partial_p13_5(39) <= partial_p17_6(39);
partial_p13_6(39) <= partial_p17_7(39);
partial_p13_7(39) <= partial_p17_8(39);
partial_p13_8(39) <= partial_p17_9(39);
partial_p13_9(39) <= partial_p17_10(39);
partial_p13_10(39) <= partial_p17_11(39);
partial_p13_11(39) <= partial_p17_12(39);
partial_p13_12(39) <= partial_p17_13(39);
FA_38 : FA port map(A=>partial_p17_0(40), B=>partial_p17_1(40), Cin => partial_p17_2(40), S=>partial_p13_2(40), Cout=>partial_p13_0(41));
HA_10 : HA port map(A=>partial_p17_3(40), B=>partial_p17_4(40), S=>partial_p13_3(40), C=>partial_p13_1(41));
partial_p13_4(40) <= partial_p17_5(40);
partial_p13_5(40) <= partial_p17_6(40);
partial_p13_6(40) <= partial_p17_7(40);
partial_p13_7(40) <= partial_p17_8(40);
partial_p13_8(40) <= partial_p17_9(40);
partial_p13_9(40) <= partial_p17_10(40);
partial_p13_10(40) <= partial_p17_11(40);
partial_p13_11(40) <= partial_p17_12(40);
partial_p13_12(40) <= partial_p17_13(40);
FA_39 : FA port map(A=>partial_p17_0(41), B=>partial_p17_1(41), Cin => partial_p17_2(41), S=>partial_p13_2(41), Cout=>partial_p13_0(42));
partial_p13_3(41) <= partial_p17_3(41);
partial_p13_4(41) <= partial_p17_4(41);
partial_p13_5(41) <= partial_p17_5(41);
partial_p13_6(41) <= partial_p17_6(41);
partial_p13_7(41) <= partial_p17_7(41);
partial_p13_8(41) <= partial_p17_8(41);
partial_p13_9(41) <= partial_p17_9(41);
partial_p13_10(41) <= partial_p17_10(41);
partial_p13_11(41) <= partial_p17_11(41);
partial_p13_12(41) <= partial_p17_12(41);
HA_11 : HA port map(A=>partial_p17_0(42), B=>partial_p17_1(42), S=>partial_p13_1(42), C=>partial_p13_0(43));
partial_p13_2(42) <= partial_p17_2(42);
partial_p13_3(42) <= partial_p17_3(42);
partial_p13_4(42) <= partial_p17_4(42);
partial_p13_5(42) <= partial_p17_5(42);
partial_p13_6(42) <= partial_p17_6(42);
partial_p13_7(42) <= partial_p17_7(42);
partial_p13_8(42) <= partial_p17_8(42);
partial_p13_9(42) <= partial_p17_9(42);
partial_p13_10(42) <= partial_p17_10(42);
partial_p13_11(42) <= partial_p17_11(42);
partial_p13_12(42) <= partial_p17_12(42);
partial_p13_1(43) <= partial_p17_0(43);
partial_p13_2(43) <= partial_p17_1(43);
partial_p13_3(43) <= partial_p17_2(43);
partial_p13_4(43) <= partial_p17_3(43);
partial_p13_5(43) <= partial_p17_4(43);
partial_p13_6(43) <= partial_p17_5(43);
partial_p13_7(43) <= partial_p17_6(43);
partial_p13_8(43) <= partial_p17_7(43);
partial_p13_9(43) <= partial_p17_8(43);
partial_p13_10(43) <= partial_p17_9(43);
partial_p13_11(43) <= partial_p17_10(43);
partial_p13_12(43) <= partial_p17_11(43);
partial_p13_0(44) <= partial_p17_0(44);
partial_p13_1(44) <= partial_p17_1(44);
partial_p13_2(44) <= partial_p17_2(44);
partial_p13_3(44) <= partial_p17_3(44);
partial_p13_4(44) <= partial_p17_4(44);
partial_p13_5(44) <= partial_p17_5(44);
partial_p13_6(44) <= partial_p17_6(44);
partial_p13_7(44) <= partial_p17_7(44);
partial_p13_8(44) <= partial_p17_8(44);
partial_p13_9(44) <= partial_p17_9(44);
partial_p13_10(44) <= partial_p17_10(44);
partial_p13_11(44) <= partial_p17_11(44);
partial_p13_12(44) <= partial_p17_12(44);
partial_p13_0(45) <= partial_p17_0(45);
partial_p13_1(45) <= partial_p17_1(45);
partial_p13_2(45) <= partial_p17_2(45);
partial_p13_3(45) <= partial_p17_3(45);
partial_p13_4(45) <= partial_p17_4(45);
partial_p13_5(45) <= partial_p17_5(45);
partial_p13_6(45) <= partial_p17_6(45);
partial_p13_7(45) <= partial_p17_7(45);
partial_p13_8(45) <= partial_p17_8(45);
partial_p13_9(45) <= partial_p17_9(45);
partial_p13_10(45) <= partial_p17_10(45);
partial_p13_11(45) <= partial_p17_11(45);
partial_p13_12(45) <= partial_p17_12(45);
partial_p13_0(46) <= partial_p17_0(46);
partial_p13_1(46) <= partial_p17_1(46);
partial_p13_2(46) <= partial_p17_2(46);
partial_p13_3(46) <= partial_p17_3(46);
partial_p13_4(46) <= partial_p17_4(46);
partial_p13_5(46) <= partial_p17_5(46);
partial_p13_6(46) <= partial_p17_6(46);
partial_p13_7(46) <= partial_p17_7(46);
partial_p13_8(46) <= partial_p17_8(46);
partial_p13_9(46) <= partial_p17_9(46);
partial_p13_10(46) <= partial_p17_10(46);
partial_p13_11(46) <= partial_p17_11(46);
partial_p13_12(46) <= partial_p17_12(46);
partial_p13_0(47) <= partial_p17_0(47);
partial_p13_1(47) <= partial_p17_1(47);
partial_p13_2(47) <= partial_p17_2(47);
partial_p13_3(47) <= partial_p17_3(47);
partial_p13_4(47) <= partial_p17_4(47);
partial_p13_5(47) <= partial_p17_5(47);
partial_p13_6(47) <= partial_p17_6(47);
partial_p13_7(47) <= partial_p17_7(47);
partial_p13_8(47) <= partial_p17_8(47);
partial_p13_9(47) <= partial_p17_9(47);
partial_p13_10(47) <= partial_p17_10(47);
partial_p13_11(47) <= partial_p17_11(47);
partial_p13_12(47) <= partial_p17_12(47);
partial_p13_0(48) <= partial_p17_0(48);
partial_p13_1(48) <= partial_p17_1(48);
partial_p13_2(48) <= partial_p17_2(48);
partial_p13_3(48) <= partial_p17_3(48);
partial_p13_4(48) <= partial_p17_4(48);
partial_p13_5(48) <= partial_p17_5(48);
partial_p13_6(48) <= partial_p17_6(48);
partial_p13_7(48) <= partial_p17_7(48);
partial_p13_8(48) <= partial_p17_8(48);
partial_p13_9(48) <= partial_p17_9(48);
partial_p13_10(48) <= partial_p17_10(48);
partial_p13_11(48) <= partial_p17_11(48);
partial_p13_12(48) <= partial_p17_12(48);
partial_p13_0(49) <= partial_p17_0(49);
partial_p13_1(49) <= partial_p17_1(49);
partial_p13_2(49) <= partial_p17_2(49);
partial_p13_3(49) <= partial_p17_3(49);
partial_p13_4(49) <= partial_p17_4(49);
partial_p13_5(49) <= partial_p17_5(49);
partial_p13_6(49) <= partial_p17_6(49);
partial_p13_7(49) <= partial_p17_7(49);
partial_p13_8(49) <= partial_p17_8(49);
partial_p13_9(49) <= partial_p17_9(49);
partial_p13_10(49) <= partial_p17_10(49);
partial_p13_11(49) <= partial_p17_11(49);
partial_p13_12(49) <= partial_p17_12(49);
partial_p13_0(50) <= partial_p17_0(50);
partial_p13_1(50) <= partial_p17_1(50);
partial_p13_2(50) <= partial_p17_2(50);
partial_p13_3(50) <= partial_p17_3(50);
partial_p13_4(50) <= partial_p17_4(50);
partial_p13_5(50) <= partial_p17_5(50);
partial_p13_6(50) <= partial_p17_6(50);
partial_p13_7(50) <= partial_p17_7(50);
partial_p13_8(50) <= partial_p17_8(50);
partial_p13_9(50) <= partial_p17_9(50);
partial_p13_10(50) <= partial_p17_10(50);
partial_p13_11(50) <= partial_p17_11(50);
partial_p13_12(50) <= partial_p17_12(50);
partial_p13_0(51) <= partial_p17_0(51);
partial_p13_1(51) <= partial_p17_1(51);
partial_p13_2(51) <= partial_p17_2(51);
partial_p13_3(51) <= partial_p17_3(51);
partial_p13_4(51) <= partial_p17_4(51);
partial_p13_5(51) <= partial_p17_5(51);
partial_p13_6(51) <= partial_p17_6(51);
partial_p13_7(51) <= partial_p17_7(51);
partial_p13_8(51) <= partial_p17_8(51);
partial_p13_9(51) <= partial_p17_9(51);
partial_p13_10(51) <= partial_p17_10(51);
partial_p13_11(51) <= partial_p17_11(51);
partial_p13_12(51) <= partial_p17_12(51);
partial_p13_0(52) <= partial_p17_0(52);
partial_p13_1(52) <= partial_p17_1(52);
partial_p13_2(52) <= partial_p17_2(52);
partial_p13_3(52) <= partial_p17_3(52);
partial_p13_4(52) <= partial_p17_4(52);
partial_p13_5(52) <= partial_p17_5(52);
partial_p13_6(52) <= partial_p17_6(52);
partial_p13_7(52) <= partial_p17_7(52);
partial_p13_8(52) <= partial_p17_8(52);
partial_p13_9(52) <= partial_p17_9(52);
partial_p13_10(52) <= partial_p17_10(52);
partial_p13_11(52) <= partial_p17_11(52);
partial_p13_12(52) <= partial_p17_12(52);
partial_p13_0(53) <= partial_p17_0(53);
partial_p13_1(53) <= partial_p17_1(53);
partial_p13_2(53) <= partial_p17_2(53);
partial_p13_3(53) <= partial_p17_3(53);
partial_p13_4(53) <= partial_p17_4(53);
partial_p13_5(53) <= partial_p17_5(53);
partial_p13_6(53) <= partial_p17_6(53);
partial_p13_7(53) <= partial_p17_7(53);
partial_p13_8(53) <= partial_p17_8(53);
partial_p13_9(53) <= partial_p17_9(53);
partial_p13_10(53) <= partial_p17_10(53);
partial_p13_11(53) <= partial_p17_11(53);
partial_p13_12(53) <= partial_p17_12(53);
partial_p13_0(54) <= partial_p17_0(54);
partial_p13_1(54) <= partial_p17_1(54);
partial_p13_2(54) <= partial_p17_2(54);
partial_p13_3(54) <= partial_p17_3(54);
partial_p13_4(54) <= partial_p17_4(54);
partial_p13_5(54) <= partial_p17_5(54);
partial_p13_6(54) <= partial_p17_6(54);
partial_p13_7(54) <= partial_p17_7(54);
partial_p13_8(54) <= partial_p17_8(54);
partial_p13_9(54) <= partial_p17_9(54);
partial_p13_10(54) <= partial_p17_10(54);
partial_p13_11(54) <= partial_p17_11(54);
partial_p13_12(54) <= partial_p17_12(54);
partial_p13_0(55) <= partial_p17_0(55);
partial_p13_1(55) <= partial_p17_1(55);
partial_p13_2(55) <= partial_p17_2(55);
partial_p13_3(55) <= partial_p17_3(55);
partial_p13_4(55) <= partial_p17_4(55);
partial_p13_5(55) <= partial_p17_5(55);
partial_p13_6(55) <= partial_p17_6(55);
partial_p13_7(55) <= partial_p17_7(55);
partial_p13_8(55) <= partial_p17_8(55);
partial_p13_9(55) <= partial_p17_9(55);
partial_p13_10(55) <= partial_p17_10(55);
partial_p13_11(55) <= partial_p17_11(55);
partial_p13_12(55) <= partial_p17_12(55);
partial_p13_0(56) <= partial_p17_0(56);
partial_p13_1(56) <= partial_p17_1(56);
partial_p13_2(56) <= partial_p17_2(56);
partial_p13_3(56) <= partial_p17_3(56);
partial_p13_4(56) <= partial_p17_4(56);
partial_p13_5(56) <= partial_p17_5(56);
partial_p13_6(56) <= partial_p17_6(56);
partial_p13_7(56) <= partial_p17_7(56);
partial_p13_8(56) <= partial_p17_8(56);
partial_p13_9(56) <= partial_p17_9(56);
partial_p13_10(56) <= partial_p17_10(56);
partial_p13_11(56) <= partial_p17_11(56);
partial_p13_12(56) <= partial_p17_12(56);
partial_p13_0(57) <= partial_p17_0(57);
partial_p13_1(57) <= partial_p17_1(57);
partial_p13_2(57) <= partial_p17_2(57);
partial_p13_3(57) <= partial_p17_3(57);
partial_p13_4(57) <= partial_p17_4(57);
partial_p13_5(57) <= partial_p17_5(57);
partial_p13_6(57) <= partial_p17_6(57);
partial_p13_7(57) <= partial_p17_7(57);
partial_p13_8(57) <= partial_p17_8(57);
partial_p13_9(57) <= partial_p17_9(57);
partial_p13_10(57) <= partial_p17_10(57);
partial_p13_11(57) <= partial_p17_11(57);
partial_p13_12(57) <= partial_p17_12(57);
partial_p13_0(58) <= partial_p17_0(58);
partial_p13_1(58) <= partial_p17_1(58);
partial_p13_2(58) <= partial_p17_2(58);
partial_p13_3(58) <= partial_p17_3(58);
partial_p13_4(58) <= partial_p17_4(58);
partial_p13_5(58) <= partial_p17_5(58);
partial_p13_6(58) <= partial_p17_6(58);
partial_p13_7(58) <= partial_p17_7(58);
partial_p13_8(58) <= partial_p17_8(58);
partial_p13_9(58) <= partial_p17_9(58);
partial_p13_10(58) <= partial_p17_10(58);
partial_p13_11(58) <= partial_p17_11(58);
partial_p13_12(58) <= partial_p17_12(58);
partial_p13_0(59) <= partial_p17_0(59);
partial_p13_1(59) <= partial_p17_1(59);
partial_p13_2(59) <= partial_p17_2(59);
partial_p13_3(59) <= partial_p17_3(59);
partial_p13_4(59) <= partial_p17_4(59);
partial_p13_5(59) <= partial_p17_5(59);
partial_p13_6(59) <= partial_p17_6(59);
partial_p13_7(59) <= partial_p17_7(59);
partial_p13_8(59) <= partial_p17_8(59);
partial_p13_9(59) <= partial_p17_9(59);
partial_p13_10(59) <= partial_p17_10(59);
partial_p13_11(59) <= partial_p17_11(59);
partial_p13_12(59) <= partial_p17_12(59);
partial_p13_0(60) <= partial_p17_0(60);
partial_p13_1(60) <= partial_p17_1(60);
partial_p13_2(60) <= partial_p17_2(60);
partial_p13_3(60) <= partial_p17_3(60);
partial_p13_4(60) <= partial_p17_4(60);
partial_p13_5(60) <= partial_p17_5(60);
partial_p13_6(60) <= partial_p17_6(60);
partial_p13_7(60) <= partial_p17_7(60);
partial_p13_8(60) <= partial_p17_8(60);
partial_p13_9(60) <= partial_p17_9(60);
partial_p13_10(60) <= partial_p17_10(60);
partial_p13_11(60) <= partial_p17_11(60);
partial_p13_12(60) <= partial_p17_12(60);
partial_p13_0(61) <= partial_p17_0(61);
partial_p13_1(61) <= partial_p17_1(61);
partial_p13_2(61) <= partial_p17_2(61);
partial_p13_3(61) <= partial_p17_3(61);
partial_p13_4(61) <= partial_p17_4(61);
partial_p13_5(61) <= partial_p17_5(61);
partial_p13_6(61) <= partial_p17_6(61);
partial_p13_7(61) <= partial_p17_7(61);
partial_p13_8(61) <= partial_p17_8(61);
partial_p13_9(61) <= partial_p17_9(61);
partial_p13_10(61) <= partial_p17_10(61);
partial_p13_11(61) <= partial_p17_11(61);
partial_p13_12(61) <= partial_p17_12(61);
partial_p13_0(62) <= partial_p17_0(62);
partial_p13_1(62) <= partial_p17_1(62);
partial_p13_2(62) <= partial_p17_2(62);
partial_p13_3(62) <= partial_p17_3(62);
partial_p13_4(62) <= partial_p17_4(62);
partial_p13_5(62) <= partial_p17_5(62);
partial_p13_6(62) <= partial_p17_6(62);
partial_p13_7(62) <= partial_p17_7(62);
partial_p13_8(62) <= partial_p17_8(62);
partial_p13_9(62) <= partial_p17_9(62);
partial_p13_10(62) <= partial_p17_10(62);
partial_p13_11(62) <= partial_p17_11(62);
partial_p13_12(62) <= partial_p17_12(62);
partial_p13_0(63) <= partial_p17_0(63);
partial_p13_1(63) <= partial_p17_1(63);
partial_p13_2(63) <= partial_p17_2(63);
partial_p13_3(63) <= partial_p17_3(63);
partial_p13_4(63) <= partial_p17_4(63);
partial_p13_5(63) <= partial_p17_5(63);
partial_p13_6(63) <= partial_p17_6(63);
partial_p13_7(63) <= partial_p17_7(63);
partial_p13_8(63) <= partial_p17_8(63);
partial_p13_9(63) <= partial_p17_9(63);
partial_p13_10(63) <= partial_p17_10(63);
partial_p13_11(63) <= partial_p17_11(63);
partial_p13_12(63) <= partial_p17_12(63);

--LEVEL 2

partial_p9_0(0) <= partial_p13_0(0);
partial_p9_1(0) <= partial_p13_1(0);
partial_p9_2(0) <= partial_p13_2(0);
partial_p9_3(0) <= partial_p13_3(0);
partial_p9_4(0) <= partial_p13_4(0);
partial_p9_5(0) <= partial_p13_5(0);
partial_p9_6(0) <= partial_p13_6(0);
partial_p9_7(0) <= partial_p13_7(0);
partial_p9_8(0) <= partial_p13_8(0);
partial_p9_0(1) <= partial_p13_0(1);
partial_p9_1(1) <= partial_p13_1(1);
partial_p9_2(1) <= partial_p13_2(1);
partial_p9_3(1) <= partial_p13_3(1);
partial_p9_4(1) <= partial_p13_4(1);
partial_p9_5(1) <= partial_p13_5(1);
partial_p9_6(1) <= partial_p13_6(1);
partial_p9_7(1) <= partial_p13_7(1);
partial_p9_8(1) <= partial_p13_8(1);
partial_p9_0(2) <= partial_p13_0(2);
partial_p9_1(2) <= partial_p13_1(2);
partial_p9_2(2) <= partial_p13_2(2);
partial_p9_3(2) <= partial_p13_3(2);
partial_p9_4(2) <= partial_p13_4(2);
partial_p9_5(2) <= partial_p13_5(2);
partial_p9_6(2) <= partial_p13_6(2);
partial_p9_7(2) <= partial_p13_7(2);
partial_p9_8(2) <= partial_p13_8(2);
partial_p9_0(3) <= partial_p13_0(3);
partial_p9_1(3) <= partial_p13_1(3);
partial_p9_2(3) <= partial_p13_2(3);
partial_p9_3(3) <= partial_p13_3(3);
partial_p9_4(3) <= partial_p13_4(3);
partial_p9_5(3) <= partial_p13_5(3);
partial_p9_6(3) <= partial_p13_6(3);
partial_p9_7(3) <= partial_p13_7(3);
partial_p9_8(3) <= partial_p13_8(3);
partial_p9_0(4) <= partial_p13_0(4);
partial_p9_1(4) <= partial_p13_1(4);
partial_p9_2(4) <= partial_p13_2(4);
partial_p9_3(4) <= partial_p13_3(4);
partial_p9_4(4) <= partial_p13_4(4);
partial_p9_5(4) <= partial_p13_5(4);
partial_p9_6(4) <= partial_p13_6(4);
partial_p9_7(4) <= partial_p13_7(4);
partial_p9_8(4) <= partial_p13_8(4);
partial_p9_0(5) <= partial_p13_0(5);
partial_p9_1(5) <= partial_p13_1(5);
partial_p9_2(5) <= partial_p13_2(5);
partial_p9_3(5) <= partial_p13_3(5);
partial_p9_4(5) <= partial_p13_4(5);
partial_p9_5(5) <= partial_p13_5(5);
partial_p9_6(5) <= partial_p13_6(5);
partial_p9_7(5) <= partial_p13_7(5);
partial_p9_8(5) <= partial_p13_8(5);
partial_p9_0(6) <= partial_p13_0(6);
partial_p9_1(6) <= partial_p13_1(6);
partial_p9_2(6) <= partial_p13_2(6);
partial_p9_3(6) <= partial_p13_3(6);
partial_p9_4(6) <= partial_p13_4(6);
partial_p9_5(6) <= partial_p13_5(6);
partial_p9_6(6) <= partial_p13_6(6);
partial_p9_7(6) <= partial_p13_7(6);
partial_p9_8(6) <= partial_p13_8(6);
partial_p9_0(7) <= partial_p13_0(7);
partial_p9_1(7) <= partial_p13_1(7);
partial_p9_2(7) <= partial_p13_2(7);
partial_p9_3(7) <= partial_p13_3(7);
partial_p9_4(7) <= partial_p13_4(7);
partial_p9_5(7) <= partial_p13_5(7);
partial_p9_6(7) <= partial_p13_6(7);
partial_p9_7(7) <= partial_p13_7(7);
partial_p9_8(7) <= partial_p13_8(7);
partial_p9_0(8) <= partial_p13_0(8);
partial_p9_1(8) <= partial_p13_1(8);
partial_p9_2(8) <= partial_p13_2(8);
partial_p9_3(8) <= partial_p13_3(8);
partial_p9_4(8) <= partial_p13_4(8);
partial_p9_5(8) <= partial_p13_5(8);
partial_p9_6(8) <= partial_p13_6(8);
partial_p9_7(8) <= partial_p13_7(8);
partial_p9_8(8) <= partial_p13_8(8);
partial_p9_0(9) <= partial_p13_0(9);
partial_p9_1(9) <= partial_p13_1(9);
partial_p9_2(9) <= partial_p13_2(9);
partial_p9_3(9) <= partial_p13_3(9);
partial_p9_4(9) <= partial_p13_4(9);
partial_p9_5(9) <= partial_p13_5(9);
partial_p9_6(9) <= partial_p13_6(9);
partial_p9_7(9) <= partial_p13_7(9);
partial_p9_8(9) <= partial_p13_8(9);
partial_p9_0(10) <= partial_p13_0(10);
partial_p9_1(10) <= partial_p13_1(10);
partial_p9_2(10) <= partial_p13_2(10);
partial_p9_3(10) <= partial_p13_3(10);
partial_p9_4(10) <= partial_p13_4(10);
partial_p9_5(10) <= partial_p13_5(10);
partial_p9_6(10) <= partial_p13_6(10);
partial_p9_7(10) <= partial_p13_7(10);
partial_p9_8(10) <= partial_p13_8(10);
partial_p9_0(11) <= partial_p13_0(11);
partial_p9_1(11) <= partial_p13_1(11);
partial_p9_2(11) <= partial_p13_2(11);
partial_p9_3(11) <= partial_p13_3(11);
partial_p9_4(11) <= partial_p13_4(11);
partial_p9_5(11) <= partial_p13_5(11);
partial_p9_6(11) <= partial_p13_6(11);
partial_p9_7(11) <= partial_p13_7(11);
partial_p9_8(11) <= partial_p13_8(11);
partial_p9_0(12) <= partial_p13_0(12);
partial_p9_1(12) <= partial_p13_1(12);
partial_p9_2(12) <= partial_p13_2(12);
partial_p9_3(12) <= partial_p13_3(12);
partial_p9_4(12) <= partial_p13_4(12);
partial_p9_5(12) <= partial_p13_5(12);
partial_p9_6(12) <= partial_p13_6(12);
partial_p9_7(12) <= partial_p13_7(12);
partial_p9_8(12) <= partial_p13_8(12);
partial_p9_0(13) <= partial_p13_0(13);
partial_p9_1(13) <= partial_p13_1(13);
partial_p9_2(13) <= partial_p13_2(13);
partial_p9_3(13) <= partial_p13_3(13);
partial_p9_4(13) <= partial_p13_4(13);
partial_p9_5(13) <= partial_p13_5(13);
partial_p9_6(13) <= partial_p13_6(13);
partial_p9_7(13) <= partial_p13_7(13);
partial_p9_8(13) <= partial_p13_8(13);
partial_p9_0(14) <= partial_p13_0(14);
partial_p9_1(14) <= partial_p13_1(14);
partial_p9_2(14) <= partial_p13_2(14);
partial_p9_3(14) <= partial_p13_3(14);
partial_p9_4(14) <= partial_p13_4(14);
partial_p9_5(14) <= partial_p13_5(14);
partial_p9_6(14) <= partial_p13_6(14);
partial_p9_7(14) <= partial_p13_7(14);
partial_p9_8(14) <= partial_p13_8(14);
partial_p9_0(15) <= partial_p13_0(15);
partial_p9_1(15) <= partial_p13_1(15);
partial_p9_2(15) <= partial_p13_2(15);
partial_p9_3(15) <= partial_p13_3(15);
partial_p9_4(15) <= partial_p13_4(15);
partial_p9_5(15) <= partial_p13_5(15);
partial_p9_6(15) <= partial_p13_6(15);
partial_p9_7(15) <= partial_p13_7(15);
partial_p9_8(15) <= partial_p13_8(15);
HA_12 : HA port map(A=>partial_p13_0(16), B=>partial_p13_1(16), S=>partial_p9_0(16), C=>partial_p9_0(17));
partial_p9_1(16) <= partial_p13_2(16);
partial_p9_2(16) <= partial_p13_3(16);
partial_p9_3(16) <= partial_p13_4(16);
partial_p9_4(16) <= partial_p13_5(16);
partial_p9_5(16) <= partial_p13_6(16);
partial_p9_6(16) <= partial_p13_7(16);
partial_p9_7(16) <= partial_p13_8(16);
partial_p9_8(16) <= partial_p13_9(16);
HA_13 : HA port map(A=>partial_p13_0(17), B=>partial_p13_1(17), S=>partial_p9_1(17), C=>partial_p9_0(18));
partial_p9_2(17) <= partial_p13_2(17);
partial_p9_3(17) <= partial_p13_3(17);
partial_p9_4(17) <= partial_p13_4(17);
partial_p9_5(17) <= partial_p13_5(17);
partial_p9_6(17) <= partial_p13_6(17);
partial_p9_7(17) <= partial_p13_7(17);
partial_p9_8(17) <= partial_p13_8(17);
FA_40 : FA port map(A=>partial_p13_0(18), B=>partial_p13_1(18), Cin => partial_p13_2(18), S=>partial_p9_1(18), Cout=>partial_p9_0(19));
HA_14 : HA port map(A=>partial_p13_3(18), B=>partial_p13_4(18), S=>partial_p9_2(18), C=>partial_p9_1(19));
partial_p9_3(18) <= partial_p13_5(18);
partial_p9_4(18) <= partial_p13_6(18);
partial_p9_5(18) <= partial_p13_7(18);
partial_p9_6(18) <= partial_p13_8(18);
partial_p9_7(18) <= partial_p13_9(18);
partial_p9_8(18) <= partial_p13_10(18);
FA_41 : FA port map(A=>partial_p13_0(19), B=>partial_p13_1(19), Cin => partial_p13_2(19), S=>partial_p9_2(19), Cout=>partial_p9_0(20));
HA_15 : HA port map(A=>partial_p13_3(19), B=>partial_p13_4(19), S=>partial_p9_3(19), C=>partial_p9_1(20));
partial_p9_4(19) <= partial_p13_5(19);
partial_p9_5(19) <= partial_p13_6(19);
partial_p9_6(19) <= partial_p13_7(19);
partial_p9_7(19) <= partial_p13_8(19);
partial_p9_8(19) <= partial_p13_9(19);
FA_42 : FA port map(A=>partial_p13_0(20), B=>partial_p13_1(20), Cin => partial_p13_2(20), S=>partial_p9_2(20), Cout=>partial_p9_0(21));
FA_43 : FA port map(A=>partial_p13_3(20), B=>partial_p13_4(20), Cin => partial_p13_5(20), S=>partial_p9_3(20), Cout=>partial_p9_1(21));
HA_16 : HA port map(A=>partial_p13_6(20), B=>partial_p13_7(20), S=>partial_p9_4(20), C=>partial_p9_2(21));
partial_p9_5(20) <= partial_p13_8(20);
partial_p9_6(20) <= partial_p13_9(20);
partial_p9_7(20) <= partial_p13_10(20);
partial_p9_8(20) <= partial_p13_11(20);
FA_44 : FA port map(A=>partial_p13_0(21), B=>partial_p13_1(21), Cin => partial_p13_2(21), S=>partial_p9_3(21), Cout=>partial_p9_0(22));
FA_45 : FA port map(A=>partial_p13_3(21), B=>partial_p13_4(21), Cin => partial_p13_5(21), S=>partial_p9_4(21), Cout=>partial_p9_1(22));
HA_17 : HA port map(A=>partial_p13_6(21), B=>partial_p13_7(21), S=>partial_p9_5(21), C=>partial_p9_2(22));
partial_p9_6(21) <= partial_p13_8(21);
partial_p9_7(21) <= partial_p13_9(21);
partial_p9_8(21) <= partial_p13_10(21);
FA_46 : FA port map(A=>partial_p13_0(22), B=>partial_p13_1(22), Cin => partial_p13_2(22), S=>partial_p9_3(22), Cout=>partial_p9_0(23));
FA_47 : FA port map(A=>partial_p13_3(22), B=>partial_p13_4(22), Cin => partial_p13_5(22), S=>partial_p9_4(22), Cout=>partial_p9_1(23));
FA_48 : FA port map(A=>partial_p13_6(22), B=>partial_p13_7(22), Cin => partial_p13_8(22), S=>partial_p9_5(22), Cout=>partial_p9_2(23));
HA_18 : HA port map(A=>partial_p13_9(22), B=>partial_p13_10(22), S=>partial_p9_6(22), C=>partial_p9_3(23));
partial_p9_7(22) <= partial_p13_11(22);
partial_p9_8(22) <= partial_p13_12(22);
FA_49 : FA port map(A=>partial_p13_0(23), B=>partial_p13_1(23), Cin => partial_p13_2(23), S=>partial_p9_4(23), Cout=>partial_p9_0(24));
FA_50 : FA port map(A=>partial_p13_3(23), B=>partial_p13_4(23), Cin => partial_p13_5(23), S=>partial_p9_5(23), Cout=>partial_p9_1(24));
FA_51 : FA port map(A=>partial_p13_6(23), B=>partial_p13_7(23), Cin => partial_p13_8(23), S=>partial_p9_6(23), Cout=>partial_p9_2(24));
HA_19 : HA port map(A=>partial_p13_9(23), B=>partial_p13_10(23), S=>partial_p9_7(23), C=>partial_p9_3(24));
partial_p9_8(23) <= partial_p13_11(23);
FA_52 : FA port map(A=>partial_p13_0(24), B=>partial_p13_1(24), Cin => partial_p13_2(24), S=>partial_p9_4(24), Cout=>partial_p9_0(25));
FA_53 : FA port map(A=>partial_p13_3(24), B=>partial_p13_4(24), Cin => partial_p13_5(24), S=>partial_p9_5(24), Cout=>partial_p9_1(25));
FA_54 : FA port map(A=>partial_p13_6(24), B=>partial_p13_7(24), Cin => partial_p13_8(24), S=>partial_p9_6(24), Cout=>partial_p9_2(25));
FA_55 : FA port map(A=>partial_p13_9(24), B=>partial_p13_10(24), Cin => partial_p13_11(24), S=>partial_p9_7(24), Cout=>partial_p9_3(25));
partial_p9_8(24) <= partial_p13_12(24);
FA_56 : FA port map(A=>partial_p13_0(25), B=>partial_p13_1(25), Cin => partial_p13_2(25), S=>partial_p9_4(25), Cout=>partial_p9_0(26));
FA_57 : FA port map(A=>partial_p13_3(25), B=>partial_p13_4(25), Cin => partial_p13_5(25), S=>partial_p9_5(25), Cout=>partial_p9_1(26));
FA_58 : FA port map(A=>partial_p13_6(25), B=>partial_p13_7(25), Cin => partial_p13_8(25), S=>partial_p9_6(25), Cout=>partial_p9_2(26));
FA_59 : FA port map(A=>partial_p13_9(25), B=>partial_p13_10(25), Cin => partial_p13_11(25), S=>partial_p9_7(25), Cout=>partial_p9_3(26));
partial_p9_8(25) <= partial_p13_12(25);
FA_60 : FA port map(A=>partial_p13_0(26), B=>partial_p13_1(26), Cin => partial_p13_2(26), S=>partial_p9_4(26), Cout=>partial_p9_0(27));
FA_61 : FA port map(A=>partial_p13_3(26), B=>partial_p13_4(26), Cin => partial_p13_5(26), S=>partial_p9_5(26), Cout=>partial_p9_1(27));
FA_62 : FA port map(A=>partial_p13_6(26), B=>partial_p13_7(26), Cin => partial_p13_8(26), S=>partial_p9_6(26), Cout=>partial_p9_2(27));
FA_63 : FA port map(A=>partial_p13_9(26), B=>partial_p13_10(26), Cin => partial_p13_11(26), S=>partial_p9_7(26), Cout=>partial_p9_3(27));
partial_p9_8(26) <= partial_p13_12(26);
FA_64 : FA port map(A=>partial_p13_0(27), B=>partial_p13_1(27), Cin => partial_p13_2(27), S=>partial_p9_4(27), Cout=>partial_p9_0(28));
FA_65 : FA port map(A=>partial_p13_3(27), B=>partial_p13_4(27), Cin => partial_p13_5(27), S=>partial_p9_5(27), Cout=>partial_p9_1(28));
FA_66 : FA port map(A=>partial_p13_6(27), B=>partial_p13_7(27), Cin => partial_p13_8(27), S=>partial_p9_6(27), Cout=>partial_p9_2(28));
FA_67 : FA port map(A=>partial_p13_9(27), B=>partial_p13_10(27), Cin => partial_p13_11(27), S=>partial_p9_7(27), Cout=>partial_p9_3(28));
partial_p9_8(27) <= partial_p13_12(27);
FA_68 : FA port map(A=>partial_p13_0(28), B=>partial_p13_1(28), Cin => partial_p13_2(28), S=>partial_p9_4(28), Cout=>partial_p9_0(29));
FA_69 : FA port map(A=>partial_p13_3(28), B=>partial_p13_4(28), Cin => partial_p13_5(28), S=>partial_p9_5(28), Cout=>partial_p9_1(29));
FA_70 : FA port map(A=>partial_p13_6(28), B=>partial_p13_7(28), Cin => partial_p13_8(28), S=>partial_p9_6(28), Cout=>partial_p9_2(29));
FA_71 : FA port map(A=>partial_p13_9(28), B=>partial_p13_10(28), Cin => partial_p13_11(28), S=>partial_p9_7(28), Cout=>partial_p9_3(29));
partial_p9_8(28) <= partial_p13_12(28);
FA_72 : FA port map(A=>partial_p13_0(29), B=>partial_p13_1(29), Cin => partial_p13_2(29), S=>partial_p9_4(29), Cout=>partial_p9_0(30));
FA_73 : FA port map(A=>partial_p13_3(29), B=>partial_p13_4(29), Cin => partial_p13_5(29), S=>partial_p9_5(29), Cout=>partial_p9_1(30));
FA_74 : FA port map(A=>partial_p13_6(29), B=>partial_p13_7(29), Cin => partial_p13_8(29), S=>partial_p9_6(29), Cout=>partial_p9_2(30));
FA_75 : FA port map(A=>partial_p13_9(29), B=>partial_p13_10(29), Cin => partial_p13_11(29), S=>partial_p9_7(29), Cout=>partial_p9_3(30));
partial_p9_8(29) <= partial_p13_12(29);
FA_76 : FA port map(A=>partial_p13_0(30), B=>partial_p13_1(30), Cin => partial_p13_2(30), S=>partial_p9_4(30), Cout=>partial_p9_0(31));
FA_77 : FA port map(A=>partial_p13_3(30), B=>partial_p13_4(30), Cin => partial_p13_5(30), S=>partial_p9_5(30), Cout=>partial_p9_1(31));
FA_78 : FA port map(A=>partial_p13_6(30), B=>partial_p13_7(30), Cin => partial_p13_8(30), S=>partial_p9_6(30), Cout=>partial_p9_2(31));
FA_79 : FA port map(A=>partial_p13_9(30), B=>partial_p13_10(30), Cin => partial_p13_11(30), S=>partial_p9_7(30), Cout=>partial_p9_3(31));
partial_p9_8(30) <= partial_p13_12(30);
FA_80 : FA port map(A=>partial_p13_0(31), B=>partial_p13_1(31), Cin => partial_p13_2(31), S=>partial_p9_4(31), Cout=>partial_p9_0(32));
FA_81 : FA port map(A=>partial_p13_3(31), B=>partial_p13_4(31), Cin => partial_p13_5(31), S=>partial_p9_5(31), Cout=>partial_p9_1(32));
FA_82 : FA port map(A=>partial_p13_6(31), B=>partial_p13_7(31), Cin => partial_p13_8(31), S=>partial_p9_6(31), Cout=>partial_p9_2(32));
FA_83 : FA port map(A=>partial_p13_9(31), B=>partial_p13_10(31), Cin => partial_p13_11(31), S=>partial_p9_7(31), Cout=>partial_p9_3(32));
partial_p9_8(31) <= partial_p13_12(31);
FA_84 : FA port map(A=>partial_p13_0(32), B=>partial_p13_1(32), Cin => partial_p13_2(32), S=>partial_p9_4(32), Cout=>partial_p9_0(33));
FA_85 : FA port map(A=>partial_p13_3(32), B=>partial_p13_4(32), Cin => partial_p13_5(32), S=>partial_p9_5(32), Cout=>partial_p9_1(33));
FA_86 : FA port map(A=>partial_p13_6(32), B=>partial_p13_7(32), Cin => partial_p13_8(32), S=>partial_p9_6(32), Cout=>partial_p9_2(33));
FA_87 : FA port map(A=>partial_p13_9(32), B=>partial_p13_10(32), Cin => partial_p13_11(32), S=>partial_p9_7(32), Cout=>partial_p9_3(33));
partial_p9_8(32) <= partial_p13_12(32);
FA_88 : FA port map(A=>partial_p13_0(33), B=>partial_p13_1(33), Cin => partial_p13_2(33), S=>partial_p9_4(33), Cout=>partial_p9_0(34));
FA_89 : FA port map(A=>partial_p13_3(33), B=>partial_p13_4(33), Cin => partial_p13_5(33), S=>partial_p9_5(33), Cout=>partial_p9_1(34));
FA_90 : FA port map(A=>partial_p13_6(33), B=>partial_p13_7(33), Cin => partial_p13_8(33), S=>partial_p9_6(33), Cout=>partial_p9_2(34));
FA_91 : FA port map(A=>partial_p13_9(33), B=>partial_p13_10(33), Cin => partial_p13_11(33), S=>partial_p9_7(33), Cout=>partial_p9_3(34));
partial_p9_8(33) <= partial_p13_12(33);
FA_92 : FA port map(A=>partial_p13_0(34), B=>partial_p13_1(34), Cin => partial_p13_2(34), S=>partial_p9_4(34), Cout=>partial_p9_0(35));
FA_93 : FA port map(A=>partial_p13_3(34), B=>partial_p13_4(34), Cin => partial_p13_5(34), S=>partial_p9_5(34), Cout=>partial_p9_1(35));
FA_94 : FA port map(A=>partial_p13_6(34), B=>partial_p13_7(34), Cin => partial_p13_8(34), S=>partial_p9_6(34), Cout=>partial_p9_2(35));
FA_95 : FA port map(A=>partial_p13_9(34), B=>partial_p13_10(34), Cin => partial_p13_11(34), S=>partial_p9_7(34), Cout=>partial_p9_3(35));
partial_p9_8(34) <= partial_p13_12(34);
FA_96 : FA port map(A=>partial_p13_0(35), B=>partial_p13_1(35), Cin => partial_p13_2(35), S=>partial_p9_4(35), Cout=>partial_p9_0(36));
FA_97 : FA port map(A=>partial_p13_3(35), B=>partial_p13_4(35), Cin => partial_p13_5(35), S=>partial_p9_5(35), Cout=>partial_p9_1(36));
FA_98 : FA port map(A=>partial_p13_6(35), B=>partial_p13_7(35), Cin => partial_p13_8(35), S=>partial_p9_6(35), Cout=>partial_p9_2(36));
FA_99 : FA port map(A=>partial_p13_9(35), B=>partial_p13_10(35), Cin => partial_p13_11(35), S=>partial_p9_7(35), Cout=>partial_p9_3(36));
partial_p9_8(35) <= partial_p13_12(35);
FA_100 : FA port map(A=>partial_p13_0(36), B=>partial_p13_1(36), Cin => partial_p13_2(36), S=>partial_p9_4(36), Cout=>partial_p9_0(37));
FA_101 : FA port map(A=>partial_p13_3(36), B=>partial_p13_4(36), Cin => partial_p13_5(36), S=>partial_p9_5(36), Cout=>partial_p9_1(37));
FA_102 : FA port map(A=>partial_p13_6(36), B=>partial_p13_7(36), Cin => partial_p13_8(36), S=>partial_p9_6(36), Cout=>partial_p9_2(37));
FA_103 : FA port map(A=>partial_p13_9(36), B=>partial_p13_10(36), Cin => partial_p13_11(36), S=>partial_p9_7(36), Cout=>partial_p9_3(37));
partial_p9_8(36) <= partial_p13_12(36);
FA_104 : FA port map(A=>partial_p13_0(37), B=>partial_p13_1(37), Cin => partial_p13_2(37), S=>partial_p9_4(37), Cout=>partial_p9_0(38));
FA_105 : FA port map(A=>partial_p13_3(37), B=>partial_p13_4(37), Cin => partial_p13_5(37), S=>partial_p9_5(37), Cout=>partial_p9_1(38));
FA_106 : FA port map(A=>partial_p13_6(37), B=>partial_p13_7(37), Cin => partial_p13_8(37), S=>partial_p9_6(37), Cout=>partial_p9_2(38));
FA_107 : FA port map(A=>partial_p13_9(37), B=>partial_p13_10(37), Cin => partial_p13_11(37), S=>partial_p9_7(37), Cout=>partial_p9_3(38));
partial_p9_8(37) <= partial_p13_12(37);
FA_108 : FA port map(A=>partial_p13_0(38), B=>partial_p13_1(38), Cin => partial_p13_2(38), S=>partial_p9_4(38), Cout=>partial_p9_0(39));
FA_109 : FA port map(A=>partial_p13_3(38), B=>partial_p13_4(38), Cin => partial_p13_5(38), S=>partial_p9_5(38), Cout=>partial_p9_1(39));
FA_110 : FA port map(A=>partial_p13_6(38), B=>partial_p13_7(38), Cin => partial_p13_8(38), S=>partial_p9_6(38), Cout=>partial_p9_2(39));
FA_111 : FA port map(A=>partial_p13_9(38), B=>partial_p13_10(38), Cin => partial_p13_11(38), S=>partial_p9_7(38), Cout=>partial_p9_3(39));
partial_p9_8(38) <= partial_p13_12(38);
FA_112 : FA port map(A=>partial_p13_0(39), B=>partial_p13_1(39), Cin => partial_p13_2(39), S=>partial_p9_4(39), Cout=>partial_p9_0(40));
FA_113 : FA port map(A=>partial_p13_3(39), B=>partial_p13_4(39), Cin => partial_p13_5(39), S=>partial_p9_5(39), Cout=>partial_p9_1(40));
FA_114 : FA port map(A=>partial_p13_6(39), B=>partial_p13_7(39), Cin => partial_p13_8(39), S=>partial_p9_6(39), Cout=>partial_p9_2(40));
FA_115 : FA port map(A=>partial_p13_9(39), B=>partial_p13_10(39), Cin => partial_p13_11(39), S=>partial_p9_7(39), Cout=>partial_p9_3(40));
partial_p9_8(39) <= partial_p13_12(39);
FA_116 : FA port map(A=>partial_p13_0(40), B=>partial_p13_1(40), Cin => partial_p13_2(40), S=>partial_p9_4(40), Cout=>partial_p9_0(41));
FA_117 : FA port map(A=>partial_p13_3(40), B=>partial_p13_4(40), Cin => partial_p13_5(40), S=>partial_p9_5(40), Cout=>partial_p9_1(41));
FA_118 : FA port map(A=>partial_p13_6(40), B=>partial_p13_7(40), Cin => partial_p13_8(40), S=>partial_p9_6(40), Cout=>partial_p9_2(41));
FA_119 : FA port map(A=>partial_p13_9(40), B=>partial_p13_10(40), Cin => partial_p13_11(40), S=>partial_p9_7(40), Cout=>partial_p9_3(41));
partial_p9_8(40) <= partial_p13_12(40);
FA_120 : FA port map(A=>partial_p13_0(41), B=>partial_p13_1(41), Cin => partial_p13_2(41), S=>partial_p9_4(41), Cout=>partial_p9_0(42));
FA_121 : FA port map(A=>partial_p13_3(41), B=>partial_p13_4(41), Cin => partial_p13_5(41), S=>partial_p9_5(41), Cout=>partial_p9_1(42));
FA_122 : FA port map(A=>partial_p13_6(41), B=>partial_p13_7(41), Cin => partial_p13_8(41), S=>partial_p9_6(41), Cout=>partial_p9_2(42));
FA_123 : FA port map(A=>partial_p13_9(41), B=>partial_p13_10(41), Cin => partial_p13_11(41), S=>partial_p9_7(41), Cout=>partial_p9_3(42));
partial_p9_8(41) <= partial_p13_12(41);
FA_124 : FA port map(A=>partial_p13_0(42), B=>partial_p13_1(42), Cin => partial_p13_2(42), S=>partial_p9_4(42), Cout=>partial_p9_0(43));
FA_125 : FA port map(A=>partial_p13_3(42), B=>partial_p13_4(42), Cin => partial_p13_5(42), S=>partial_p9_5(42), Cout=>partial_p9_1(43));
FA_126 : FA port map(A=>partial_p13_6(42), B=>partial_p13_7(42), Cin => partial_p13_8(42), S=>partial_p9_6(42), Cout=>partial_p9_2(43));
FA_127 : FA port map(A=>partial_p13_9(42), B=>partial_p13_10(42), Cin => partial_p13_11(42), S=>partial_p9_7(42), Cout=>partial_p9_3(43));
partial_p9_8(42) <= partial_p13_12(42);
FA_128 : FA port map(A=>partial_p13_0(43), B=>partial_p13_1(43), Cin => partial_p13_2(43), S=>partial_p9_4(43), Cout=>partial_p9_0(44));
FA_129 : FA port map(A=>partial_p13_3(43), B=>partial_p13_4(43), Cin => partial_p13_5(43), S=>partial_p9_5(43), Cout=>partial_p9_1(44));
FA_130 : FA port map(A=>partial_p13_6(43), B=>partial_p13_7(43), Cin => partial_p13_8(43), S=>partial_p9_6(43), Cout=>partial_p9_2(44));
FA_131 : FA port map(A=>partial_p13_9(43), B=>partial_p13_10(43), Cin => partial_p13_11(43), S=>partial_p9_7(43), Cout=>partial_p9_3(44));
partial_p9_8(43) <= partial_p13_12(43);
FA_132 : FA port map(A=>partial_p13_0(44), B=>partial_p13_1(44), Cin => partial_p13_2(44), S=>partial_p9_4(44), Cout=>partial_p9_0(45));
FA_133 : FA port map(A=>partial_p13_3(44), B=>partial_p13_4(44), Cin => partial_p13_5(44), S=>partial_p9_5(44), Cout=>partial_p9_1(45));
FA_134 : FA port map(A=>partial_p13_6(44), B=>partial_p13_7(44), Cin => partial_p13_8(44), S=>partial_p9_6(44), Cout=>partial_p9_2(45));
HA_20 : HA port map(A=>partial_p13_9(44), B=>partial_p13_10(44), S=>partial_p9_7(44), C=>partial_p9_3(45));
partial_p9_8(44) <= partial_p13_11(44);
FA_135 : FA port map(A=>partial_p13_0(45), B=>partial_p13_1(45), Cin => partial_p13_2(45), S=>partial_p9_4(45), Cout=>partial_p9_0(46));
FA_136 : FA port map(A=>partial_p13_3(45), B=>partial_p13_4(45), Cin => partial_p13_5(45), S=>partial_p9_5(45), Cout=>partial_p9_1(46));
FA_137 : FA port map(A=>partial_p13_6(45), B=>partial_p13_7(45), Cin => partial_p13_8(45), S=>partial_p9_6(45), Cout=>partial_p9_2(46));
partial_p9_7(45) <= partial_p13_9(45);
partial_p9_8(45) <= partial_p13_10(45);
FA_138 : FA port map(A=>partial_p13_0(46), B=>partial_p13_1(46), Cin => partial_p13_2(46), S=>partial_p9_3(46), Cout=>partial_p9_0(47));
FA_139 : FA port map(A=>partial_p13_3(46), B=>partial_p13_4(46), Cin => partial_p13_5(46), S=>partial_p9_4(46), Cout=>partial_p9_1(47));
HA_21 : HA port map(A=>partial_p13_6(46), B=>partial_p13_7(46), S=>partial_p9_5(46), C=>partial_p9_2(47));
partial_p9_6(46) <= partial_p13_8(46);
partial_p9_7(46) <= partial_p13_9(46);
partial_p9_8(46) <= partial_p13_10(46);
FA_140 : FA port map(A=>partial_p13_0(47), B=>partial_p13_1(47), Cin => partial_p13_2(47), S=>partial_p9_3(47), Cout=>partial_p9_0(48));
FA_141 : FA port map(A=>partial_p13_3(47), B=>partial_p13_4(47), Cin => partial_p13_5(47), S=>partial_p9_4(47), Cout=>partial_p9_1(48));
partial_p9_5(47) <= partial_p13_6(47);
partial_p9_6(47) <= partial_p13_7(47);
partial_p9_7(47) <= partial_p13_8(47);
partial_p9_8(47) <= partial_p13_9(47);
FA_142 : FA port map(A=>partial_p13_0(48), B=>partial_p13_1(48), Cin => partial_p13_2(48), S=>partial_p9_2(48), Cout=>partial_p9_0(49));
HA_22 : HA port map(A=>partial_p13_3(48), B=>partial_p13_4(48), S=>partial_p9_3(48), C=>partial_p9_1(49));
partial_p9_4(48) <= partial_p13_5(48);
partial_p9_5(48) <= partial_p13_6(48);
partial_p9_6(48) <= partial_p13_7(48);
partial_p9_7(48) <= partial_p13_8(48);
partial_p9_8(48) <= partial_p13_9(48);
FA_143 : FA port map(A=>partial_p13_0(49), B=>partial_p13_1(49), Cin => partial_p13_2(49), S=>partial_p9_2(49), Cout=>partial_p9_0(50));
partial_p9_3(49) <= partial_p13_3(49);
partial_p9_4(49) <= partial_p13_4(49);
partial_p9_5(49) <= partial_p13_5(49);
partial_p9_6(49) <= partial_p13_6(49);
partial_p9_7(49) <= partial_p13_7(49);
partial_p9_8(49) <= partial_p13_8(49);
HA_23 : HA port map(A=>partial_p13_0(50), B=>partial_p13_1(50), S=>partial_p9_1(50), C=>partial_p9_0(51));
partial_p9_2(50) <= partial_p13_2(50);
partial_p9_3(50) <= partial_p13_3(50);
partial_p9_4(50) <= partial_p13_4(50);
partial_p9_5(50) <= partial_p13_5(50);
partial_p9_6(50) <= partial_p13_6(50);
partial_p9_7(50) <= partial_p13_7(50);
partial_p9_8(50) <= partial_p13_8(50);
partial_p9_1(51) <= partial_p13_0(51);
partial_p9_2(51) <= partial_p13_1(51);
partial_p9_3(51) <= partial_p13_2(51);
partial_p9_4(51) <= partial_p13_3(51);
partial_p9_5(51) <= partial_p13_4(51);
partial_p9_6(51) <= partial_p13_5(51);
partial_p9_7(51) <= partial_p13_6(51);
partial_p9_8(51) <= partial_p13_7(51);
partial_p9_0(52) <= partial_p13_0(52);
partial_p9_1(52) <= partial_p13_1(52);
partial_p9_2(52) <= partial_p13_2(52);
partial_p9_3(52) <= partial_p13_3(52);
partial_p9_4(52) <= partial_p13_4(52);
partial_p9_5(52) <= partial_p13_5(52);
partial_p9_6(52) <= partial_p13_6(52);
partial_p9_7(52) <= partial_p13_7(52);
partial_p9_8(52) <= partial_p13_8(52);
partial_p9_0(53) <= partial_p13_0(53);
partial_p9_1(53) <= partial_p13_1(53);
partial_p9_2(53) <= partial_p13_2(53);
partial_p9_3(53) <= partial_p13_3(53);
partial_p9_4(53) <= partial_p13_4(53);
partial_p9_5(53) <= partial_p13_5(53);
partial_p9_6(53) <= partial_p13_6(53);
partial_p9_7(53) <= partial_p13_7(53);
partial_p9_8(53) <= partial_p13_8(53);
partial_p9_0(54) <= partial_p13_0(54);
partial_p9_1(54) <= partial_p13_1(54);
partial_p9_2(54) <= partial_p13_2(54);
partial_p9_3(54) <= partial_p13_3(54);
partial_p9_4(54) <= partial_p13_4(54);
partial_p9_5(54) <= partial_p13_5(54);
partial_p9_6(54) <= partial_p13_6(54);
partial_p9_7(54) <= partial_p13_7(54);
partial_p9_8(54) <= partial_p13_8(54);
partial_p9_0(55) <= partial_p13_0(55);
partial_p9_1(55) <= partial_p13_1(55);
partial_p9_2(55) <= partial_p13_2(55);
partial_p9_3(55) <= partial_p13_3(55);
partial_p9_4(55) <= partial_p13_4(55);
partial_p9_5(55) <= partial_p13_5(55);
partial_p9_6(55) <= partial_p13_6(55);
partial_p9_7(55) <= partial_p13_7(55);
partial_p9_8(55) <= partial_p13_8(55);
partial_p9_0(56) <= partial_p13_0(56);
partial_p9_1(56) <= partial_p13_1(56);
partial_p9_2(56) <= partial_p13_2(56);
partial_p9_3(56) <= partial_p13_3(56);
partial_p9_4(56) <= partial_p13_4(56);
partial_p9_5(56) <= partial_p13_5(56);
partial_p9_6(56) <= partial_p13_6(56);
partial_p9_7(56) <= partial_p13_7(56);
partial_p9_8(56) <= partial_p13_8(56);
partial_p9_0(57) <= partial_p13_0(57);
partial_p9_1(57) <= partial_p13_1(57);
partial_p9_2(57) <= partial_p13_2(57);
partial_p9_3(57) <= partial_p13_3(57);
partial_p9_4(57) <= partial_p13_4(57);
partial_p9_5(57) <= partial_p13_5(57);
partial_p9_6(57) <= partial_p13_6(57);
partial_p9_7(57) <= partial_p13_7(57);
partial_p9_8(57) <= partial_p13_8(57);
partial_p9_0(58) <= partial_p13_0(58);
partial_p9_1(58) <= partial_p13_1(58);
partial_p9_2(58) <= partial_p13_2(58);
partial_p9_3(58) <= partial_p13_3(58);
partial_p9_4(58) <= partial_p13_4(58);
partial_p9_5(58) <= partial_p13_5(58);
partial_p9_6(58) <= partial_p13_6(58);
partial_p9_7(58) <= partial_p13_7(58);
partial_p9_8(58) <= partial_p13_8(58);
partial_p9_0(59) <= partial_p13_0(59);
partial_p9_1(59) <= partial_p13_1(59);
partial_p9_2(59) <= partial_p13_2(59);
partial_p9_3(59) <= partial_p13_3(59);
partial_p9_4(59) <= partial_p13_4(59);
partial_p9_5(59) <= partial_p13_5(59);
partial_p9_6(59) <= partial_p13_6(59);
partial_p9_7(59) <= partial_p13_7(59);
partial_p9_8(59) <= partial_p13_8(59);
partial_p9_0(60) <= partial_p13_0(60);
partial_p9_1(60) <= partial_p13_1(60);
partial_p9_2(60) <= partial_p13_2(60);
partial_p9_3(60) <= partial_p13_3(60);
partial_p9_4(60) <= partial_p13_4(60);
partial_p9_5(60) <= partial_p13_5(60);
partial_p9_6(60) <= partial_p13_6(60);
partial_p9_7(60) <= partial_p13_7(60);
partial_p9_8(60) <= partial_p13_8(60);
partial_p9_0(61) <= partial_p13_0(61);
partial_p9_1(61) <= partial_p13_1(61);
partial_p9_2(61) <= partial_p13_2(61);
partial_p9_3(61) <= partial_p13_3(61);
partial_p9_4(61) <= partial_p13_4(61);
partial_p9_5(61) <= partial_p13_5(61);
partial_p9_6(61) <= partial_p13_6(61);
partial_p9_7(61) <= partial_p13_7(61);
partial_p9_8(61) <= partial_p13_8(61);
partial_p9_0(62) <= partial_p13_0(62);
partial_p9_1(62) <= partial_p13_1(62);
partial_p9_2(62) <= partial_p13_2(62);
partial_p9_3(62) <= partial_p13_3(62);
partial_p9_4(62) <= partial_p13_4(62);
partial_p9_5(62) <= partial_p13_5(62);
partial_p9_6(62) <= partial_p13_6(62);
partial_p9_7(62) <= partial_p13_7(62);
partial_p9_8(62) <= partial_p13_8(62);
partial_p9_0(63) <= partial_p13_0(63);
partial_p9_1(63) <= partial_p13_1(63);
partial_p9_2(63) <= partial_p13_2(63);
partial_p9_3(63) <= partial_p13_3(63);
partial_p9_4(63) <= partial_p13_4(63);
partial_p9_5(63) <= partial_p13_5(63);
partial_p9_6(63) <= partial_p13_6(63);
partial_p9_7(63) <= partial_p13_7(63);
partial_p9_8(63) <= partial_p13_8(63);

--LEVEL 3

partial_p6_0(0) <= partial_p9_0(0);
partial_p6_1(0) <= partial_p9_1(0);
partial_p6_2(0) <= partial_p9_2(0);
partial_p6_3(0) <= partial_p9_3(0);
partial_p6_4(0) <= partial_p9_4(0);
partial_p6_5(0) <= partial_p9_5(0);
partial_p6_0(1) <= partial_p9_0(1);
partial_p6_1(1) <= partial_p9_1(1);
partial_p6_2(1) <= partial_p9_2(1);
partial_p6_3(1) <= partial_p9_3(1);
partial_p6_4(1) <= partial_p9_4(1);
partial_p6_5(1) <= partial_p9_5(1);
partial_p6_0(2) <= partial_p9_0(2);
partial_p6_1(2) <= partial_p9_1(2);
partial_p6_2(2) <= partial_p9_2(2);
partial_p6_3(2) <= partial_p9_3(2);
partial_p6_4(2) <= partial_p9_4(2);
partial_p6_5(2) <= partial_p9_5(2);
partial_p6_0(3) <= partial_p9_0(3);
partial_p6_1(3) <= partial_p9_1(3);
partial_p6_2(3) <= partial_p9_2(3);
partial_p6_3(3) <= partial_p9_3(3);
partial_p6_4(3) <= partial_p9_4(3);
partial_p6_5(3) <= partial_p9_5(3);
partial_p6_0(4) <= partial_p9_0(4);
partial_p6_1(4) <= partial_p9_1(4);
partial_p6_2(4) <= partial_p9_2(4);
partial_p6_3(4) <= partial_p9_3(4);
partial_p6_4(4) <= partial_p9_4(4);
partial_p6_5(4) <= partial_p9_5(4);
partial_p6_0(5) <= partial_p9_0(5);
partial_p6_1(5) <= partial_p9_1(5);
partial_p6_2(5) <= partial_p9_2(5);
partial_p6_3(5) <= partial_p9_3(5);
partial_p6_4(5) <= partial_p9_4(5);
partial_p6_5(5) <= partial_p9_5(5);
partial_p6_0(6) <= partial_p9_0(6);
partial_p6_1(6) <= partial_p9_1(6);
partial_p6_2(6) <= partial_p9_2(6);
partial_p6_3(6) <= partial_p9_3(6);
partial_p6_4(6) <= partial_p9_4(6);
partial_p6_5(6) <= partial_p9_5(6);
partial_p6_0(7) <= partial_p9_0(7);
partial_p6_1(7) <= partial_p9_1(7);
partial_p6_2(7) <= partial_p9_2(7);
partial_p6_3(7) <= partial_p9_3(7);
partial_p6_4(7) <= partial_p9_4(7);
partial_p6_5(7) <= partial_p9_5(7);
partial_p6_0(8) <= partial_p9_0(8);
partial_p6_1(8) <= partial_p9_1(8);
partial_p6_2(8) <= partial_p9_2(8);
partial_p6_3(8) <= partial_p9_3(8);
partial_p6_4(8) <= partial_p9_4(8);
partial_p6_5(8) <= partial_p9_5(8);
partial_p6_0(9) <= partial_p9_0(9);
partial_p6_1(9) <= partial_p9_1(9);
partial_p6_2(9) <= partial_p9_2(9);
partial_p6_3(9) <= partial_p9_3(9);
partial_p6_4(9) <= partial_p9_4(9);
partial_p6_5(9) <= partial_p9_5(9);
HA_24 : HA port map(A=>partial_p9_0(10), B=>partial_p9_1(10), S=>partial_p6_0(10), C=>partial_p6_0(11));
partial_p6_1(10) <= partial_p9_2(10);
partial_p6_2(10) <= partial_p9_3(10);
partial_p6_3(10) <= partial_p9_4(10);
partial_p6_4(10) <= partial_p9_5(10);
partial_p6_5(10) <= partial_p9_6(10);
HA_25 : HA port map(A=>partial_p9_0(11), B=>partial_p9_1(11), S=>partial_p6_1(11), C=>partial_p6_0(12));
partial_p6_2(11) <= partial_p9_2(11);
partial_p6_3(11) <= partial_p9_3(11);
partial_p6_4(11) <= partial_p9_4(11);
partial_p6_5(11) <= partial_p9_5(11);
FA_144 : FA port map(A=>partial_p9_0(12), B=>partial_p9_1(12), Cin => partial_p9_2(12), S=>partial_p6_1(12), Cout=>partial_p6_0(13));
HA_26 : HA port map(A=>partial_p9_3(12), B=>partial_p9_4(12), S=>partial_p6_2(12), C=>partial_p6_1(13));
partial_p6_3(12) <= partial_p9_5(12);
partial_p6_4(12) <= partial_p9_6(12);
partial_p6_5(12) <= partial_p9_7(12);
FA_145 : FA port map(A=>partial_p9_0(13), B=>partial_p9_1(13), Cin => partial_p9_2(13), S=>partial_p6_2(13), Cout=>partial_p6_0(14));
HA_27 : HA port map(A=>partial_p9_3(13), B=>partial_p9_4(13), S=>partial_p6_3(13), C=>partial_p6_1(14));
partial_p6_4(13) <= partial_p9_5(13);
partial_p6_5(13) <= partial_p9_6(13);
FA_146 : FA port map(A=>partial_p9_0(14), B=>partial_p9_1(14), Cin => partial_p9_2(14), S=>partial_p6_2(14), Cout=>partial_p6_0(15));
FA_147 : FA port map(A=>partial_p9_3(14), B=>partial_p9_4(14), Cin => partial_p9_5(14), S=>partial_p6_3(14), Cout=>partial_p6_1(15));
HA_28 : HA port map(A=>partial_p9_6(14), B=>partial_p9_7(14), S=>partial_p6_4(14), C=>partial_p6_2(15));
partial_p6_5(14) <= partial_p9_8(14);
FA_148 : FA port map(A=>partial_p9_0(15), B=>partial_p9_1(15), Cin => partial_p9_2(15), S=>partial_p6_3(15), Cout=>partial_p6_0(16));
FA_149 : FA port map(A=>partial_p9_3(15), B=>partial_p9_4(15), Cin => partial_p9_5(15), S=>partial_p6_4(15), Cout=>partial_p6_1(16));
HA_29 : HA port map(A=>partial_p9_6(15), B=>partial_p9_7(15), S=>partial_p6_5(15), C=>partial_p6_2(16));
FA_150 : FA port map(A=>partial_p9_0(16), B=>partial_p9_1(16), Cin => partial_p9_2(16), S=>partial_p6_3(16), Cout=>partial_p6_0(17));
FA_151 : FA port map(A=>partial_p9_3(16), B=>partial_p9_4(16), Cin => partial_p9_5(16), S=>partial_p6_4(16), Cout=>partial_p6_1(17));
FA_152 : FA port map(A=>partial_p9_6(16), B=>partial_p9_7(16), Cin => partial_p9_8(16), S=>partial_p6_5(16), Cout=>partial_p6_2(17));
FA_153 : FA port map(A=>partial_p9_0(17), B=>partial_p9_1(17), Cin => partial_p9_2(17), S=>partial_p6_3(17), Cout=>partial_p6_0(18));
FA_154 : FA port map(A=>partial_p9_3(17), B=>partial_p9_4(17), Cin => partial_p9_5(17), S=>partial_p6_4(17), Cout=>partial_p6_1(18));
FA_155 : FA port map(A=>partial_p9_6(17), B=>partial_p9_7(17), Cin => partial_p9_8(17), S=>partial_p6_5(17), Cout=>partial_p6_2(18));
FA_156 : FA port map(A=>partial_p9_0(18), B=>partial_p9_1(18), Cin => partial_p9_2(18), S=>partial_p6_3(18), Cout=>partial_p6_0(19));
FA_157 : FA port map(A=>partial_p9_3(18), B=>partial_p9_4(18), Cin => partial_p9_5(18), S=>partial_p6_4(18), Cout=>partial_p6_1(19));
FA_158 : FA port map(A=>partial_p9_6(18), B=>partial_p9_7(18), Cin => partial_p9_8(18), S=>partial_p6_5(18), Cout=>partial_p6_2(19));
FA_159 : FA port map(A=>partial_p9_0(19), B=>partial_p9_1(19), Cin => partial_p9_2(19), S=>partial_p6_3(19), Cout=>partial_p6_0(20));
FA_160 : FA port map(A=>partial_p9_3(19), B=>partial_p9_4(19), Cin => partial_p9_5(19), S=>partial_p6_4(19), Cout=>partial_p6_1(20));
FA_161 : FA port map(A=>partial_p9_6(19), B=>partial_p9_7(19), Cin => partial_p9_8(19), S=>partial_p6_5(19), Cout=>partial_p6_2(20));
FA_162 : FA port map(A=>partial_p9_0(20), B=>partial_p9_1(20), Cin => partial_p9_2(20), S=>partial_p6_3(20), Cout=>partial_p6_0(21));
FA_163 : FA port map(A=>partial_p9_3(20), B=>partial_p9_4(20), Cin => partial_p9_5(20), S=>partial_p6_4(20), Cout=>partial_p6_1(21));
FA_164 : FA port map(A=>partial_p9_6(20), B=>partial_p9_7(20), Cin => partial_p9_8(20), S=>partial_p6_5(20), Cout=>partial_p6_2(21));
FA_165 : FA port map(A=>partial_p9_0(21), B=>partial_p9_1(21), Cin => partial_p9_2(21), S=>partial_p6_3(21), Cout=>partial_p6_0(22));
FA_166 : FA port map(A=>partial_p9_3(21), B=>partial_p9_4(21), Cin => partial_p9_5(21), S=>partial_p6_4(21), Cout=>partial_p6_1(22));
FA_167 : FA port map(A=>partial_p9_6(21), B=>partial_p9_7(21), Cin => partial_p9_8(21), S=>partial_p6_5(21), Cout=>partial_p6_2(22));
FA_168 : FA port map(A=>partial_p9_0(22), B=>partial_p9_1(22), Cin => partial_p9_2(22), S=>partial_p6_3(22), Cout=>partial_p6_0(23));
FA_169 : FA port map(A=>partial_p9_3(22), B=>partial_p9_4(22), Cin => partial_p9_5(22), S=>partial_p6_4(22), Cout=>partial_p6_1(23));
FA_170 : FA port map(A=>partial_p9_6(22), B=>partial_p9_7(22), Cin => partial_p9_8(22), S=>partial_p6_5(22), Cout=>partial_p6_2(23));
FA_171 : FA port map(A=>partial_p9_0(23), B=>partial_p9_1(23), Cin => partial_p9_2(23), S=>partial_p6_3(23), Cout=>partial_p6_0(24));
FA_172 : FA port map(A=>partial_p9_3(23), B=>partial_p9_4(23), Cin => partial_p9_5(23), S=>partial_p6_4(23), Cout=>partial_p6_1(24));
FA_173 : FA port map(A=>partial_p9_6(23), B=>partial_p9_7(23), Cin => partial_p9_8(23), S=>partial_p6_5(23), Cout=>partial_p6_2(24));
FA_174 : FA port map(A=>partial_p9_0(24), B=>partial_p9_1(24), Cin => partial_p9_2(24), S=>partial_p6_3(24), Cout=>partial_p6_0(25));
FA_175 : FA port map(A=>partial_p9_3(24), B=>partial_p9_4(24), Cin => partial_p9_5(24), S=>partial_p6_4(24), Cout=>partial_p6_1(25));
FA_176 : FA port map(A=>partial_p9_6(24), B=>partial_p9_7(24), Cin => partial_p9_8(24), S=>partial_p6_5(24), Cout=>partial_p6_2(25));
FA_177 : FA port map(A=>partial_p9_0(25), B=>partial_p9_1(25), Cin => partial_p9_2(25), S=>partial_p6_3(25), Cout=>partial_p6_0(26));
FA_178 : FA port map(A=>partial_p9_3(25), B=>partial_p9_4(25), Cin => partial_p9_5(25), S=>partial_p6_4(25), Cout=>partial_p6_1(26));
FA_179 : FA port map(A=>partial_p9_6(25), B=>partial_p9_7(25), Cin => partial_p9_8(25), S=>partial_p6_5(25), Cout=>partial_p6_2(26));
FA_180 : FA port map(A=>partial_p9_0(26), B=>partial_p9_1(26), Cin => partial_p9_2(26), S=>partial_p6_3(26), Cout=>partial_p6_0(27));
FA_181 : FA port map(A=>partial_p9_3(26), B=>partial_p9_4(26), Cin => partial_p9_5(26), S=>partial_p6_4(26), Cout=>partial_p6_1(27));
FA_182 : FA port map(A=>partial_p9_6(26), B=>partial_p9_7(26), Cin => partial_p9_8(26), S=>partial_p6_5(26), Cout=>partial_p6_2(27));
FA_183 : FA port map(A=>partial_p9_0(27), B=>partial_p9_1(27), Cin => partial_p9_2(27), S=>partial_p6_3(27), Cout=>partial_p6_0(28));
FA_184 : FA port map(A=>partial_p9_3(27), B=>partial_p9_4(27), Cin => partial_p9_5(27), S=>partial_p6_4(27), Cout=>partial_p6_1(28));
FA_185 : FA port map(A=>partial_p9_6(27), B=>partial_p9_7(27), Cin => partial_p9_8(27), S=>partial_p6_5(27), Cout=>partial_p6_2(28));
FA_186 : FA port map(A=>partial_p9_0(28), B=>partial_p9_1(28), Cin => partial_p9_2(28), S=>partial_p6_3(28), Cout=>partial_p6_0(29));
FA_187 : FA port map(A=>partial_p9_3(28), B=>partial_p9_4(28), Cin => partial_p9_5(28), S=>partial_p6_4(28), Cout=>partial_p6_1(29));
FA_188 : FA port map(A=>partial_p9_6(28), B=>partial_p9_7(28), Cin => partial_p9_8(28), S=>partial_p6_5(28), Cout=>partial_p6_2(29));
FA_189 : FA port map(A=>partial_p9_0(29), B=>partial_p9_1(29), Cin => partial_p9_2(29), S=>partial_p6_3(29), Cout=>partial_p6_0(30));
FA_190 : FA port map(A=>partial_p9_3(29), B=>partial_p9_4(29), Cin => partial_p9_5(29), S=>partial_p6_4(29), Cout=>partial_p6_1(30));
FA_191 : FA port map(A=>partial_p9_6(29), B=>partial_p9_7(29), Cin => partial_p9_8(29), S=>partial_p6_5(29), Cout=>partial_p6_2(30));
FA_192 : FA port map(A=>partial_p9_0(30), B=>partial_p9_1(30), Cin => partial_p9_2(30), S=>partial_p6_3(30), Cout=>partial_p6_0(31));
FA_193 : FA port map(A=>partial_p9_3(30), B=>partial_p9_4(30), Cin => partial_p9_5(30), S=>partial_p6_4(30), Cout=>partial_p6_1(31));
FA_194 : FA port map(A=>partial_p9_6(30), B=>partial_p9_7(30), Cin => partial_p9_8(30), S=>partial_p6_5(30), Cout=>partial_p6_2(31));
FA_195 : FA port map(A=>partial_p9_0(31), B=>partial_p9_1(31), Cin => partial_p9_2(31), S=>partial_p6_3(31), Cout=>partial_p6_0(32));
FA_196 : FA port map(A=>partial_p9_3(31), B=>partial_p9_4(31), Cin => partial_p9_5(31), S=>partial_p6_4(31), Cout=>partial_p6_1(32));
FA_197 : FA port map(A=>partial_p9_6(31), B=>partial_p9_7(31), Cin => partial_p9_8(31), S=>partial_p6_5(31), Cout=>partial_p6_2(32));
FA_198 : FA port map(A=>partial_p9_0(32), B=>partial_p9_1(32), Cin => partial_p9_2(32), S=>partial_p6_3(32), Cout=>partial_p6_0(33));
FA_199 : FA port map(A=>partial_p9_3(32), B=>partial_p9_4(32), Cin => partial_p9_5(32), S=>partial_p6_4(32), Cout=>partial_p6_1(33));
FA_200 : FA port map(A=>partial_p9_6(32), B=>partial_p9_7(32), Cin => partial_p9_8(32), S=>partial_p6_5(32), Cout=>partial_p6_2(33));
FA_201 : FA port map(A=>partial_p9_0(33), B=>partial_p9_1(33), Cin => partial_p9_2(33), S=>partial_p6_3(33), Cout=>partial_p6_0(34));
FA_202 : FA port map(A=>partial_p9_3(33), B=>partial_p9_4(33), Cin => partial_p9_5(33), S=>partial_p6_4(33), Cout=>partial_p6_1(34));
FA_203 : FA port map(A=>partial_p9_6(33), B=>partial_p9_7(33), Cin => partial_p9_8(33), S=>partial_p6_5(33), Cout=>partial_p6_2(34));
FA_204 : FA port map(A=>partial_p9_0(34), B=>partial_p9_1(34), Cin => partial_p9_2(34), S=>partial_p6_3(34), Cout=>partial_p6_0(35));
FA_205 : FA port map(A=>partial_p9_3(34), B=>partial_p9_4(34), Cin => partial_p9_5(34), S=>partial_p6_4(34), Cout=>partial_p6_1(35));
FA_206 : FA port map(A=>partial_p9_6(34), B=>partial_p9_7(34), Cin => partial_p9_8(34), S=>partial_p6_5(34), Cout=>partial_p6_2(35));
FA_207 : FA port map(A=>partial_p9_0(35), B=>partial_p9_1(35), Cin => partial_p9_2(35), S=>partial_p6_3(35), Cout=>partial_p6_0(36));
FA_208 : FA port map(A=>partial_p9_3(35), B=>partial_p9_4(35), Cin => partial_p9_5(35), S=>partial_p6_4(35), Cout=>partial_p6_1(36));
FA_209 : FA port map(A=>partial_p9_6(35), B=>partial_p9_7(35), Cin => partial_p9_8(35), S=>partial_p6_5(35), Cout=>partial_p6_2(36));
FA_210 : FA port map(A=>partial_p9_0(36), B=>partial_p9_1(36), Cin => partial_p9_2(36), S=>partial_p6_3(36), Cout=>partial_p6_0(37));
FA_211 : FA port map(A=>partial_p9_3(36), B=>partial_p9_4(36), Cin => partial_p9_5(36), S=>partial_p6_4(36), Cout=>partial_p6_1(37));
FA_212 : FA port map(A=>partial_p9_6(36), B=>partial_p9_7(36), Cin => partial_p9_8(36), S=>partial_p6_5(36), Cout=>partial_p6_2(37));
FA_213 : FA port map(A=>partial_p9_0(37), B=>partial_p9_1(37), Cin => partial_p9_2(37), S=>partial_p6_3(37), Cout=>partial_p6_0(38));
FA_214 : FA port map(A=>partial_p9_3(37), B=>partial_p9_4(37), Cin => partial_p9_5(37), S=>partial_p6_4(37), Cout=>partial_p6_1(38));
FA_215 : FA port map(A=>partial_p9_6(37), B=>partial_p9_7(37), Cin => partial_p9_8(37), S=>partial_p6_5(37), Cout=>partial_p6_2(38));
FA_216 : FA port map(A=>partial_p9_0(38), B=>partial_p9_1(38), Cin => partial_p9_2(38), S=>partial_p6_3(38), Cout=>partial_p6_0(39));
FA_217 : FA port map(A=>partial_p9_3(38), B=>partial_p9_4(38), Cin => partial_p9_5(38), S=>partial_p6_4(38), Cout=>partial_p6_1(39));
FA_218 : FA port map(A=>partial_p9_6(38), B=>partial_p9_7(38), Cin => partial_p9_8(38), S=>partial_p6_5(38), Cout=>partial_p6_2(39));
FA_219 : FA port map(A=>partial_p9_0(39), B=>partial_p9_1(39), Cin => partial_p9_2(39), S=>partial_p6_3(39), Cout=>partial_p6_0(40));
FA_220 : FA port map(A=>partial_p9_3(39), B=>partial_p9_4(39), Cin => partial_p9_5(39), S=>partial_p6_4(39), Cout=>partial_p6_1(40));
FA_221 : FA port map(A=>partial_p9_6(39), B=>partial_p9_7(39), Cin => partial_p9_8(39), S=>partial_p6_5(39), Cout=>partial_p6_2(40));
FA_222 : FA port map(A=>partial_p9_0(40), B=>partial_p9_1(40), Cin => partial_p9_2(40), S=>partial_p6_3(40), Cout=>partial_p6_0(41));
FA_223 : FA port map(A=>partial_p9_3(40), B=>partial_p9_4(40), Cin => partial_p9_5(40), S=>partial_p6_4(40), Cout=>partial_p6_1(41));
FA_224 : FA port map(A=>partial_p9_6(40), B=>partial_p9_7(40), Cin => partial_p9_8(40), S=>partial_p6_5(40), Cout=>partial_p6_2(41));
FA_225 : FA port map(A=>partial_p9_0(41), B=>partial_p9_1(41), Cin => partial_p9_2(41), S=>partial_p6_3(41), Cout=>partial_p6_0(42));
FA_226 : FA port map(A=>partial_p9_3(41), B=>partial_p9_4(41), Cin => partial_p9_5(41), S=>partial_p6_4(41), Cout=>partial_p6_1(42));
FA_227 : FA port map(A=>partial_p9_6(41), B=>partial_p9_7(41), Cin => partial_p9_8(41), S=>partial_p6_5(41), Cout=>partial_p6_2(42));
FA_228 : FA port map(A=>partial_p9_0(42), B=>partial_p9_1(42), Cin => partial_p9_2(42), S=>partial_p6_3(42), Cout=>partial_p6_0(43));
FA_229 : FA port map(A=>partial_p9_3(42), B=>partial_p9_4(42), Cin => partial_p9_5(42), S=>partial_p6_4(42), Cout=>partial_p6_1(43));
FA_230 : FA port map(A=>partial_p9_6(42), B=>partial_p9_7(42), Cin => partial_p9_8(42), S=>partial_p6_5(42), Cout=>partial_p6_2(43));
FA_231 : FA port map(A=>partial_p9_0(43), B=>partial_p9_1(43), Cin => partial_p9_2(43), S=>partial_p6_3(43), Cout=>partial_p6_0(44));
FA_232 : FA port map(A=>partial_p9_3(43), B=>partial_p9_4(43), Cin => partial_p9_5(43), S=>partial_p6_4(43), Cout=>partial_p6_1(44));
FA_233 : FA port map(A=>partial_p9_6(43), B=>partial_p9_7(43), Cin => partial_p9_8(43), S=>partial_p6_5(43), Cout=>partial_p6_2(44));
FA_234 : FA port map(A=>partial_p9_0(44), B=>partial_p9_1(44), Cin => partial_p9_2(44), S=>partial_p6_3(44), Cout=>partial_p6_0(45));
FA_235 : FA port map(A=>partial_p9_3(44), B=>partial_p9_4(44), Cin => partial_p9_5(44), S=>partial_p6_4(44), Cout=>partial_p6_1(45));
FA_236 : FA port map(A=>partial_p9_6(44), B=>partial_p9_7(44), Cin => partial_p9_8(44), S=>partial_p6_5(44), Cout=>partial_p6_2(45));
FA_237 : FA port map(A=>partial_p9_0(45), B=>partial_p9_1(45), Cin => partial_p9_2(45), S=>partial_p6_3(45), Cout=>partial_p6_0(46));
FA_238 : FA port map(A=>partial_p9_3(45), B=>partial_p9_4(45), Cin => partial_p9_5(45), S=>partial_p6_4(45), Cout=>partial_p6_1(46));
FA_239 : FA port map(A=>partial_p9_6(45), B=>partial_p9_7(45), Cin => partial_p9_8(45), S=>partial_p6_5(45), Cout=>partial_p6_2(46));
FA_240 : FA port map(A=>partial_p9_0(46), B=>partial_p9_1(46), Cin => partial_p9_2(46), S=>partial_p6_3(46), Cout=>partial_p6_0(47));
FA_241 : FA port map(A=>partial_p9_3(46), B=>partial_p9_4(46), Cin => partial_p9_5(46), S=>partial_p6_4(46), Cout=>partial_p6_1(47));
FA_242 : FA port map(A=>partial_p9_6(46), B=>partial_p9_7(46), Cin => partial_p9_8(46), S=>partial_p6_5(46), Cout=>partial_p6_2(47));
FA_243 : FA port map(A=>partial_p9_0(47), B=>partial_p9_1(47), Cin => partial_p9_2(47), S=>partial_p6_3(47), Cout=>partial_p6_0(48));
FA_244 : FA port map(A=>partial_p9_3(47), B=>partial_p9_4(47), Cin => partial_p9_5(47), S=>partial_p6_4(47), Cout=>partial_p6_1(48));
FA_245 : FA port map(A=>partial_p9_6(47), B=>partial_p9_7(47), Cin => partial_p9_8(47), S=>partial_p6_5(47), Cout=>partial_p6_2(48));
FA_246 : FA port map(A=>partial_p9_0(48), B=>partial_p9_1(48), Cin => partial_p9_2(48), S=>partial_p6_3(48), Cout=>partial_p6_0(49));
FA_247 : FA port map(A=>partial_p9_3(48), B=>partial_p9_4(48), Cin => partial_p9_5(48), S=>partial_p6_4(48), Cout=>partial_p6_1(49));
FA_248 : FA port map(A=>partial_p9_6(48), B=>partial_p9_7(48), Cin => partial_p9_8(48), S=>partial_p6_5(48), Cout=>partial_p6_2(49));
FA_249 : FA port map(A=>partial_p9_0(49), B=>partial_p9_1(49), Cin => partial_p9_2(49), S=>partial_p6_3(49), Cout=>partial_p6_0(50));
FA_250 : FA port map(A=>partial_p9_3(49), B=>partial_p9_4(49), Cin => partial_p9_5(49), S=>partial_p6_4(49), Cout=>partial_p6_1(50));
FA_251 : FA port map(A=>partial_p9_6(49), B=>partial_p9_7(49), Cin => partial_p9_8(49), S=>partial_p6_5(49), Cout=>partial_p6_2(50));
FA_252 : FA port map(A=>partial_p9_0(50), B=>partial_p9_1(50), Cin => partial_p9_2(50), S=>partial_p6_3(50), Cout=>partial_p6_0(51));
FA_253 : FA port map(A=>partial_p9_3(50), B=>partial_p9_4(50), Cin => partial_p9_5(50), S=>partial_p6_4(50), Cout=>partial_p6_1(51));
FA_254 : FA port map(A=>partial_p9_6(50), B=>partial_p9_7(50), Cin => partial_p9_8(50), S=>partial_p6_5(50), Cout=>partial_p6_2(51));
FA_255 : FA port map(A=>partial_p9_0(51), B=>partial_p9_1(51), Cin => partial_p9_2(51), S=>partial_p6_3(51), Cout=>partial_p6_0(52));
FA_256 : FA port map(A=>partial_p9_3(51), B=>partial_p9_4(51), Cin => partial_p9_5(51), S=>partial_p6_4(51), Cout=>partial_p6_1(52));
FA_257 : FA port map(A=>partial_p9_6(51), B=>partial_p9_7(51), Cin => partial_p9_8(51), S=>partial_p6_5(51), Cout=>partial_p6_2(52));
FA_258 : FA port map(A=>partial_p9_0(52), B=>partial_p9_1(52), Cin => partial_p9_2(52), S=>partial_p6_3(52), Cout=>partial_p6_0(53));
FA_259 : FA port map(A=>partial_p9_3(52), B=>partial_p9_4(52), Cin => partial_p9_5(52), S=>partial_p6_4(52), Cout=>partial_p6_1(53));
HA_30 : HA port map(A=>partial_p9_6(52), B=>partial_p9_7(52), S=>partial_p6_5(52), C=>partial_p6_2(53));
FA_260 : FA port map(A=>partial_p9_0(53), B=>partial_p9_1(53), Cin => partial_p9_2(53), S=>partial_p6_3(53), Cout=>partial_p6_0(54));
FA_261 : FA port map(A=>partial_p9_3(53), B=>partial_p9_4(53), Cin => partial_p9_5(53), S=>partial_p6_4(53), Cout=>partial_p6_1(54));
partial_p6_5(53) <= partial_p9_6(53);
FA_262 : FA port map(A=>partial_p9_0(54), B=>partial_p9_1(54), Cin => partial_p9_2(54), S=>partial_p6_2(54), Cout=>partial_p6_0(55));
HA_31 : HA port map(A=>partial_p9_3(54), B=>partial_p9_4(54), S=>partial_p6_3(54), C=>partial_p6_1(55));
partial_p6_4(54) <= partial_p9_5(54);
partial_p6_5(54) <= partial_p9_6(54);
FA_263 : FA port map(A=>partial_p9_0(55), B=>partial_p9_1(55), Cin => partial_p9_2(55), S=>partial_p6_2(55), Cout=>partial_p6_0(56));
partial_p6_3(55) <= partial_p9_3(55);
partial_p6_4(55) <= partial_p9_4(55);
partial_p6_5(55) <= partial_p9_5(55);
HA_32 : HA port map(A=>partial_p9_0(56), B=>partial_p9_1(56), S=>partial_p6_1(56), C=>partial_p6_0(57));
partial_p6_2(56) <= partial_p9_2(56);
partial_p6_3(56) <= partial_p9_3(56);
partial_p6_4(56) <= partial_p9_4(56);
partial_p6_5(56) <= partial_p9_5(56);
partial_p6_1(57) <= partial_p9_0(57);
partial_p6_2(57) <= partial_p9_1(57);
partial_p6_3(57) <= partial_p9_2(57);
partial_p6_4(57) <= partial_p9_3(57);
partial_p6_5(57) <= partial_p9_4(57);
partial_p6_0(58) <= partial_p9_0(58);
partial_p6_1(58) <= partial_p9_1(58);
partial_p6_2(58) <= partial_p9_2(58);
partial_p6_3(58) <= partial_p9_3(58);
partial_p6_4(58) <= partial_p9_4(58);
partial_p6_5(58) <= partial_p9_5(58);
partial_p6_0(59) <= partial_p9_0(59);
partial_p6_1(59) <= partial_p9_1(59);
partial_p6_2(59) <= partial_p9_2(59);
partial_p6_3(59) <= partial_p9_3(59);
partial_p6_4(59) <= partial_p9_4(59);
partial_p6_5(59) <= partial_p9_5(59);
partial_p6_0(60) <= partial_p9_0(60);
partial_p6_1(60) <= partial_p9_1(60);
partial_p6_2(60) <= partial_p9_2(60);
partial_p6_3(60) <= partial_p9_3(60);
partial_p6_4(60) <= partial_p9_4(60);
partial_p6_5(60) <= partial_p9_5(60);
partial_p6_0(61) <= partial_p9_0(61);
partial_p6_1(61) <= partial_p9_1(61);
partial_p6_2(61) <= partial_p9_2(61);
partial_p6_3(61) <= partial_p9_3(61);
partial_p6_4(61) <= partial_p9_4(61);
partial_p6_5(61) <= partial_p9_5(61);
partial_p6_0(62) <= partial_p9_0(62);
partial_p6_1(62) <= partial_p9_1(62);
partial_p6_2(62) <= partial_p9_2(62);
partial_p6_3(62) <= partial_p9_3(62);
partial_p6_4(62) <= partial_p9_4(62);
partial_p6_5(62) <= partial_p9_5(62);
partial_p6_0(63) <= partial_p9_0(63);
partial_p6_1(63) <= partial_p9_1(63);
partial_p6_2(63) <= partial_p9_2(63);
partial_p6_3(63) <= partial_p9_3(63);
partial_p6_4(63) <= partial_p9_4(63);
partial_p6_5(63) <= partial_p9_5(63);

--LEVEL 4

partial_p4_0(0) <= partial_p6_0(0);
partial_p4_1(0) <= partial_p6_1(0);
partial_p4_2(0) <= partial_p6_2(0);
partial_p4_3(0) <= partial_p6_3(0);
partial_p4_0(1) <= partial_p6_0(1);
partial_p4_1(1) <= partial_p6_1(1);
partial_p4_2(1) <= partial_p6_2(1);
partial_p4_3(1) <= partial_p6_3(1);
partial_p4_0(2) <= partial_p6_0(2);
partial_p4_1(2) <= partial_p6_1(2);
partial_p4_2(2) <= partial_p6_2(2);
partial_p4_3(2) <= partial_p6_3(2);
partial_p4_0(3) <= partial_p6_0(3);
partial_p4_1(3) <= partial_p6_1(3);
partial_p4_2(3) <= partial_p6_2(3);
partial_p4_3(3) <= partial_p6_3(3);
partial_p4_0(4) <= partial_p6_0(4);
partial_p4_1(4) <= partial_p6_1(4);
partial_p4_2(4) <= partial_p6_2(4);
partial_p4_3(4) <= partial_p6_3(4);
partial_p4_0(5) <= partial_p6_0(5);
partial_p4_1(5) <= partial_p6_1(5);
partial_p4_2(5) <= partial_p6_2(5);
partial_p4_3(5) <= partial_p6_3(5);
HA_33 : HA port map(A=>partial_p6_0(6), B=>partial_p6_1(6), S=>partial_p4_0(6), C=>partial_p4_0(7));
partial_p4_1(6) <= partial_p6_2(6);
partial_p4_2(6) <= partial_p6_3(6);
partial_p4_3(6) <= partial_p6_4(6);
HA_34 : HA port map(A=>partial_p6_0(7), B=>partial_p6_1(7), S=>partial_p4_1(7), C=>partial_p4_0(8));
partial_p4_2(7) <= partial_p6_2(7);
partial_p4_3(7) <= partial_p6_3(7);
FA_264 : FA port map(A=>partial_p6_0(8), B=>partial_p6_1(8), Cin => partial_p6_2(8), S=>partial_p4_1(8), Cout=>partial_p4_0(9));
HA_35 : HA port map(A=>partial_p6_3(8), B=>partial_p6_4(8), S=>partial_p4_2(8), C=>partial_p4_1(9));
partial_p4_3(8) <= partial_p6_5(8);
FA_265 : FA port map(A=>partial_p6_0(9), B=>partial_p6_1(9), Cin => partial_p6_2(9), S=>partial_p4_2(9), Cout=>partial_p4_0(10));
HA_36 : HA port map(A=>partial_p6_3(9), B=>partial_p6_4(9), S=>partial_p4_3(9), C=>partial_p4_1(10));
FA_266 : FA port map(A=>partial_p6_0(10), B=>partial_p6_1(10), Cin => partial_p6_2(10), S=>partial_p4_2(10), Cout=>partial_p4_0(11));
FA_267 : FA port map(A=>partial_p6_3(10), B=>partial_p6_4(10), Cin => partial_p6_5(10), S=>partial_p4_3(10), Cout=>partial_p4_1(11));
FA_268 : FA port map(A=>partial_p6_0(11), B=>partial_p6_1(11), Cin => partial_p6_2(11), S=>partial_p4_2(11), Cout=>partial_p4_0(12));
FA_269 : FA port map(A=>partial_p6_3(11), B=>partial_p6_4(11), Cin => partial_p6_5(11), S=>partial_p4_3(11), Cout=>partial_p4_1(12));
FA_270 : FA port map(A=>partial_p6_0(12), B=>partial_p6_1(12), Cin => partial_p6_2(12), S=>partial_p4_2(12), Cout=>partial_p4_0(13));
FA_271 : FA port map(A=>partial_p6_3(12), B=>partial_p6_4(12), Cin => partial_p6_5(12), S=>partial_p4_3(12), Cout=>partial_p4_1(13));
FA_272 : FA port map(A=>partial_p6_0(13), B=>partial_p6_1(13), Cin => partial_p6_2(13), S=>partial_p4_2(13), Cout=>partial_p4_0(14));
FA_273 : FA port map(A=>partial_p6_3(13), B=>partial_p6_4(13), Cin => partial_p6_5(13), S=>partial_p4_3(13), Cout=>partial_p4_1(14));
FA_274 : FA port map(A=>partial_p6_0(14), B=>partial_p6_1(14), Cin => partial_p6_2(14), S=>partial_p4_2(14), Cout=>partial_p4_0(15));
FA_275 : FA port map(A=>partial_p6_3(14), B=>partial_p6_4(14), Cin => partial_p6_5(14), S=>partial_p4_3(14), Cout=>partial_p4_1(15));
FA_276 : FA port map(A=>partial_p6_0(15), B=>partial_p6_1(15), Cin => partial_p6_2(15), S=>partial_p4_2(15), Cout=>partial_p4_0(16));
FA_277 : FA port map(A=>partial_p6_3(15), B=>partial_p6_4(15), Cin => partial_p6_5(15), S=>partial_p4_3(15), Cout=>partial_p4_1(16));
FA_278 : FA port map(A=>partial_p6_0(16), B=>partial_p6_1(16), Cin => partial_p6_2(16), S=>partial_p4_2(16), Cout=>partial_p4_0(17));
FA_279 : FA port map(A=>partial_p6_3(16), B=>partial_p6_4(16), Cin => partial_p6_5(16), S=>partial_p4_3(16), Cout=>partial_p4_1(17));
FA_280 : FA port map(A=>partial_p6_0(17), B=>partial_p6_1(17), Cin => partial_p6_2(17), S=>partial_p4_2(17), Cout=>partial_p4_0(18));
FA_281 : FA port map(A=>partial_p6_3(17), B=>partial_p6_4(17), Cin => partial_p6_5(17), S=>partial_p4_3(17), Cout=>partial_p4_1(18));
FA_282 : FA port map(A=>partial_p6_0(18), B=>partial_p6_1(18), Cin => partial_p6_2(18), S=>partial_p4_2(18), Cout=>partial_p4_0(19));
FA_283 : FA port map(A=>partial_p6_3(18), B=>partial_p6_4(18), Cin => partial_p6_5(18), S=>partial_p4_3(18), Cout=>partial_p4_1(19));
FA_284 : FA port map(A=>partial_p6_0(19), B=>partial_p6_1(19), Cin => partial_p6_2(19), S=>partial_p4_2(19), Cout=>partial_p4_0(20));
FA_285 : FA port map(A=>partial_p6_3(19), B=>partial_p6_4(19), Cin => partial_p6_5(19), S=>partial_p4_3(19), Cout=>partial_p4_1(20));
FA_286 : FA port map(A=>partial_p6_0(20), B=>partial_p6_1(20), Cin => partial_p6_2(20), S=>partial_p4_2(20), Cout=>partial_p4_0(21));
FA_287 : FA port map(A=>partial_p6_3(20), B=>partial_p6_4(20), Cin => partial_p6_5(20), S=>partial_p4_3(20), Cout=>partial_p4_1(21));
FA_288 : FA port map(A=>partial_p6_0(21), B=>partial_p6_1(21), Cin => partial_p6_2(21), S=>partial_p4_2(21), Cout=>partial_p4_0(22));
FA_289 : FA port map(A=>partial_p6_3(21), B=>partial_p6_4(21), Cin => partial_p6_5(21), S=>partial_p4_3(21), Cout=>partial_p4_1(22));
FA_290 : FA port map(A=>partial_p6_0(22), B=>partial_p6_1(22), Cin => partial_p6_2(22), S=>partial_p4_2(22), Cout=>partial_p4_0(23));
FA_291 : FA port map(A=>partial_p6_3(22), B=>partial_p6_4(22), Cin => partial_p6_5(22), S=>partial_p4_3(22), Cout=>partial_p4_1(23));
FA_292 : FA port map(A=>partial_p6_0(23), B=>partial_p6_1(23), Cin => partial_p6_2(23), S=>partial_p4_2(23), Cout=>partial_p4_0(24));
FA_293 : FA port map(A=>partial_p6_3(23), B=>partial_p6_4(23), Cin => partial_p6_5(23), S=>partial_p4_3(23), Cout=>partial_p4_1(24));
FA_294 : FA port map(A=>partial_p6_0(24), B=>partial_p6_1(24), Cin => partial_p6_2(24), S=>partial_p4_2(24), Cout=>partial_p4_0(25));
FA_295 : FA port map(A=>partial_p6_3(24), B=>partial_p6_4(24), Cin => partial_p6_5(24), S=>partial_p4_3(24), Cout=>partial_p4_1(25));
FA_296 : FA port map(A=>partial_p6_0(25), B=>partial_p6_1(25), Cin => partial_p6_2(25), S=>partial_p4_2(25), Cout=>partial_p4_0(26));
FA_297 : FA port map(A=>partial_p6_3(25), B=>partial_p6_4(25), Cin => partial_p6_5(25), S=>partial_p4_3(25), Cout=>partial_p4_1(26));
FA_298 : FA port map(A=>partial_p6_0(26), B=>partial_p6_1(26), Cin => partial_p6_2(26), S=>partial_p4_2(26), Cout=>partial_p4_0(27));
FA_299 : FA port map(A=>partial_p6_3(26), B=>partial_p6_4(26), Cin => partial_p6_5(26), S=>partial_p4_3(26), Cout=>partial_p4_1(27));
FA_300 : FA port map(A=>partial_p6_0(27), B=>partial_p6_1(27), Cin => partial_p6_2(27), S=>partial_p4_2(27), Cout=>partial_p4_0(28));
FA_301 : FA port map(A=>partial_p6_3(27), B=>partial_p6_4(27), Cin => partial_p6_5(27), S=>partial_p4_3(27), Cout=>partial_p4_1(28));
FA_302 : FA port map(A=>partial_p6_0(28), B=>partial_p6_1(28), Cin => partial_p6_2(28), S=>partial_p4_2(28), Cout=>partial_p4_0(29));
FA_303 : FA port map(A=>partial_p6_3(28), B=>partial_p6_4(28), Cin => partial_p6_5(28), S=>partial_p4_3(28), Cout=>partial_p4_1(29));
FA_304 : FA port map(A=>partial_p6_0(29), B=>partial_p6_1(29), Cin => partial_p6_2(29), S=>partial_p4_2(29), Cout=>partial_p4_0(30));
FA_305 : FA port map(A=>partial_p6_3(29), B=>partial_p6_4(29), Cin => partial_p6_5(29), S=>partial_p4_3(29), Cout=>partial_p4_1(30));
FA_306 : FA port map(A=>partial_p6_0(30), B=>partial_p6_1(30), Cin => partial_p6_2(30), S=>partial_p4_2(30), Cout=>partial_p4_0(31));
FA_307 : FA port map(A=>partial_p6_3(30), B=>partial_p6_4(30), Cin => partial_p6_5(30), S=>partial_p4_3(30), Cout=>partial_p4_1(31));
FA_308 : FA port map(A=>partial_p6_0(31), B=>partial_p6_1(31), Cin => partial_p6_2(31), S=>partial_p4_2(31), Cout=>partial_p4_0(32));
FA_309 : FA port map(A=>partial_p6_3(31), B=>partial_p6_4(31), Cin => partial_p6_5(31), S=>partial_p4_3(31), Cout=>partial_p4_1(32));
FA_310 : FA port map(A=>partial_p6_0(32), B=>partial_p6_1(32), Cin => partial_p6_2(32), S=>partial_p4_2(32), Cout=>partial_p4_0(33));
FA_311 : FA port map(A=>partial_p6_3(32), B=>partial_p6_4(32), Cin => partial_p6_5(32), S=>partial_p4_3(32), Cout=>partial_p4_1(33));
FA_312 : FA port map(A=>partial_p6_0(33), B=>partial_p6_1(33), Cin => partial_p6_2(33), S=>partial_p4_2(33), Cout=>partial_p4_0(34));
FA_313 : FA port map(A=>partial_p6_3(33), B=>partial_p6_4(33), Cin => partial_p6_5(33), S=>partial_p4_3(33), Cout=>partial_p4_1(34));
FA_314 : FA port map(A=>partial_p6_0(34), B=>partial_p6_1(34), Cin => partial_p6_2(34), S=>partial_p4_2(34), Cout=>partial_p4_0(35));
FA_315 : FA port map(A=>partial_p6_3(34), B=>partial_p6_4(34), Cin => partial_p6_5(34), S=>partial_p4_3(34), Cout=>partial_p4_1(35));
FA_316 : FA port map(A=>partial_p6_0(35), B=>partial_p6_1(35), Cin => partial_p6_2(35), S=>partial_p4_2(35), Cout=>partial_p4_0(36));
FA_317 : FA port map(A=>partial_p6_3(35), B=>partial_p6_4(35), Cin => partial_p6_5(35), S=>partial_p4_3(35), Cout=>partial_p4_1(36));
FA_318 : FA port map(A=>partial_p6_0(36), B=>partial_p6_1(36), Cin => partial_p6_2(36), S=>partial_p4_2(36), Cout=>partial_p4_0(37));
FA_319 : FA port map(A=>partial_p6_3(36), B=>partial_p6_4(36), Cin => partial_p6_5(36), S=>partial_p4_3(36), Cout=>partial_p4_1(37));
FA_320 : FA port map(A=>partial_p6_0(37), B=>partial_p6_1(37), Cin => partial_p6_2(37), S=>partial_p4_2(37), Cout=>partial_p4_0(38));
FA_321 : FA port map(A=>partial_p6_3(37), B=>partial_p6_4(37), Cin => partial_p6_5(37), S=>partial_p4_3(37), Cout=>partial_p4_1(38));
FA_322 : FA port map(A=>partial_p6_0(38), B=>partial_p6_1(38), Cin => partial_p6_2(38), S=>partial_p4_2(38), Cout=>partial_p4_0(39));
FA_323 : FA port map(A=>partial_p6_3(38), B=>partial_p6_4(38), Cin => partial_p6_5(38), S=>partial_p4_3(38), Cout=>partial_p4_1(39));
FA_324 : FA port map(A=>partial_p6_0(39), B=>partial_p6_1(39), Cin => partial_p6_2(39), S=>partial_p4_2(39), Cout=>partial_p4_0(40));
FA_325 : FA port map(A=>partial_p6_3(39), B=>partial_p6_4(39), Cin => partial_p6_5(39), S=>partial_p4_3(39), Cout=>partial_p4_1(40));
FA_326 : FA port map(A=>partial_p6_0(40), B=>partial_p6_1(40), Cin => partial_p6_2(40), S=>partial_p4_2(40), Cout=>partial_p4_0(41));
FA_327 : FA port map(A=>partial_p6_3(40), B=>partial_p6_4(40), Cin => partial_p6_5(40), S=>partial_p4_3(40), Cout=>partial_p4_1(41));
FA_328 : FA port map(A=>partial_p6_0(41), B=>partial_p6_1(41), Cin => partial_p6_2(41), S=>partial_p4_2(41), Cout=>partial_p4_0(42));
FA_329 : FA port map(A=>partial_p6_3(41), B=>partial_p6_4(41), Cin => partial_p6_5(41), S=>partial_p4_3(41), Cout=>partial_p4_1(42));
FA_330 : FA port map(A=>partial_p6_0(42), B=>partial_p6_1(42), Cin => partial_p6_2(42), S=>partial_p4_2(42), Cout=>partial_p4_0(43));
FA_331 : FA port map(A=>partial_p6_3(42), B=>partial_p6_4(42), Cin => partial_p6_5(42), S=>partial_p4_3(42), Cout=>partial_p4_1(43));
FA_332 : FA port map(A=>partial_p6_0(43), B=>partial_p6_1(43), Cin => partial_p6_2(43), S=>partial_p4_2(43), Cout=>partial_p4_0(44));
FA_333 : FA port map(A=>partial_p6_3(43), B=>partial_p6_4(43), Cin => partial_p6_5(43), S=>partial_p4_3(43), Cout=>partial_p4_1(44));
FA_334 : FA port map(A=>partial_p6_0(44), B=>partial_p6_1(44), Cin => partial_p6_2(44), S=>partial_p4_2(44), Cout=>partial_p4_0(45));
FA_335 : FA port map(A=>partial_p6_3(44), B=>partial_p6_4(44), Cin => partial_p6_5(44), S=>partial_p4_3(44), Cout=>partial_p4_1(45));
FA_336 : FA port map(A=>partial_p6_0(45), B=>partial_p6_1(45), Cin => partial_p6_2(45), S=>partial_p4_2(45), Cout=>partial_p4_0(46));
FA_337 : FA port map(A=>partial_p6_3(45), B=>partial_p6_4(45), Cin => partial_p6_5(45), S=>partial_p4_3(45), Cout=>partial_p4_1(46));
FA_338 : FA port map(A=>partial_p6_0(46), B=>partial_p6_1(46), Cin => partial_p6_2(46), S=>partial_p4_2(46), Cout=>partial_p4_0(47));
FA_339 : FA port map(A=>partial_p6_3(46), B=>partial_p6_4(46), Cin => partial_p6_5(46), S=>partial_p4_3(46), Cout=>partial_p4_1(47));
FA_340 : FA port map(A=>partial_p6_0(47), B=>partial_p6_1(47), Cin => partial_p6_2(47), S=>partial_p4_2(47), Cout=>partial_p4_0(48));
FA_341 : FA port map(A=>partial_p6_3(47), B=>partial_p6_4(47), Cin => partial_p6_5(47), S=>partial_p4_3(47), Cout=>partial_p4_1(48));
FA_342 : FA port map(A=>partial_p6_0(48), B=>partial_p6_1(48), Cin => partial_p6_2(48), S=>partial_p4_2(48), Cout=>partial_p4_0(49));
FA_343 : FA port map(A=>partial_p6_3(48), B=>partial_p6_4(48), Cin => partial_p6_5(48), S=>partial_p4_3(48), Cout=>partial_p4_1(49));
FA_344 : FA port map(A=>partial_p6_0(49), B=>partial_p6_1(49), Cin => partial_p6_2(49), S=>partial_p4_2(49), Cout=>partial_p4_0(50));
FA_345 : FA port map(A=>partial_p6_3(49), B=>partial_p6_4(49), Cin => partial_p6_5(49), S=>partial_p4_3(49), Cout=>partial_p4_1(50));
FA_346 : FA port map(A=>partial_p6_0(50), B=>partial_p6_1(50), Cin => partial_p6_2(50), S=>partial_p4_2(50), Cout=>partial_p4_0(51));
FA_347 : FA port map(A=>partial_p6_3(50), B=>partial_p6_4(50), Cin => partial_p6_5(50), S=>partial_p4_3(50), Cout=>partial_p4_1(51));
FA_348 : FA port map(A=>partial_p6_0(51), B=>partial_p6_1(51), Cin => partial_p6_2(51), S=>partial_p4_2(51), Cout=>partial_p4_0(52));
FA_349 : FA port map(A=>partial_p6_3(51), B=>partial_p6_4(51), Cin => partial_p6_5(51), S=>partial_p4_3(51), Cout=>partial_p4_1(52));
FA_350 : FA port map(A=>partial_p6_0(52), B=>partial_p6_1(52), Cin => partial_p6_2(52), S=>partial_p4_2(52), Cout=>partial_p4_0(53));
FA_351 : FA port map(A=>partial_p6_3(52), B=>partial_p6_4(52), Cin => partial_p6_5(52), S=>partial_p4_3(52), Cout=>partial_p4_1(53));
FA_352 : FA port map(A=>partial_p6_0(53), B=>partial_p6_1(53), Cin => partial_p6_2(53), S=>partial_p4_2(53), Cout=>partial_p4_0(54));
FA_353 : FA port map(A=>partial_p6_3(53), B=>partial_p6_4(53), Cin => partial_p6_5(53), S=>partial_p4_3(53), Cout=>partial_p4_1(54));
FA_354 : FA port map(A=>partial_p6_0(54), B=>partial_p6_1(54), Cin => partial_p6_2(54), S=>partial_p4_2(54), Cout=>partial_p4_0(55));
FA_355 : FA port map(A=>partial_p6_3(54), B=>partial_p6_4(54), Cin => partial_p6_5(54), S=>partial_p4_3(54), Cout=>partial_p4_1(55));
FA_356 : FA port map(A=>partial_p6_0(55), B=>partial_p6_1(55), Cin => partial_p6_2(55), S=>partial_p4_2(55), Cout=>partial_p4_0(56));
FA_357 : FA port map(A=>partial_p6_3(55), B=>partial_p6_4(55), Cin => partial_p6_5(55), S=>partial_p4_3(55), Cout=>partial_p4_1(56));
FA_358 : FA port map(A=>partial_p6_0(56), B=>partial_p6_1(56), Cin => partial_p6_2(56), S=>partial_p4_2(56), Cout=>partial_p4_0(57));
FA_359 : FA port map(A=>partial_p6_3(56), B=>partial_p6_4(56), Cin => partial_p6_5(56), S=>partial_p4_3(56), Cout=>partial_p4_1(57));
FA_360 : FA port map(A=>partial_p6_0(57), B=>partial_p6_1(57), Cin => partial_p6_2(57), S=>partial_p4_2(57), Cout=>partial_p4_0(58));
FA_361 : FA port map(A=>partial_p6_3(57), B=>partial_p6_4(57), Cin => partial_p6_5(57), S=>partial_p4_3(57), Cout=>partial_p4_1(58));
FA_362 : FA port map(A=>partial_p6_0(58), B=>partial_p6_1(58), Cin => partial_p6_2(58), S=>partial_p4_2(58), Cout=>partial_p4_0(59));
HA_37 : HA port map(A=>partial_p6_3(58), B=>partial_p6_4(58), S=>partial_p4_3(58), C=>partial_p4_1(59));
FA_363 : FA port map(A=>partial_p6_0(59), B=>partial_p6_1(59), Cin => partial_p6_2(59), S=>partial_p4_2(59), Cout=>partial_p4_0(60));
partial_p4_3(59) <= partial_p6_3(59);
HA_38 : HA port map(A=>partial_p6_0(60), B=>partial_p6_1(60), S=>partial_p4_1(60), C=>partial_p4_0(61));
partial_p4_2(60) <= partial_p6_2(60);
partial_p4_3(60) <= partial_p6_3(60);
partial_p4_1(61) <= partial_p6_0(61);
partial_p4_2(61) <= partial_p6_1(61);
partial_p4_3(61) <= partial_p6_2(61);
partial_p4_0(62) <= partial_p6_0(62);
partial_p4_1(62) <= partial_p6_1(62);
partial_p4_2(62) <= partial_p6_2(62);
partial_p4_3(62) <= partial_p6_3(62);
partial_p4_0(63) <= partial_p6_0(63);
partial_p4_1(63) <= partial_p6_1(63);
partial_p4_2(63) <= partial_p6_2(63);
partial_p4_3(63) <= partial_p6_3(63);

--LEVEL 5

partial_p3_0(0) <= partial_p4_0(0);
partial_p3_1(0) <= partial_p4_1(0);
partial_p3_2(0) <= partial_p4_2(0);
partial_p3_0(1) <= partial_p4_0(1);
partial_p3_1(1) <= partial_p4_1(1);
partial_p3_2(1) <= partial_p4_2(1);
partial_p3_0(2) <= partial_p4_0(2);
partial_p3_1(2) <= partial_p4_1(2);
partial_p3_2(2) <= partial_p4_2(2);
partial_p3_0(3) <= partial_p4_0(3);
partial_p3_1(3) <= partial_p4_1(3);
partial_p3_2(3) <= partial_p4_2(3);
HA_39 : HA port map(A=>partial_p4_0(4), B=>partial_p4_1(4), S=>partial_p3_0(4), C=>partial_p3_0(5));
partial_p3_1(4) <= partial_p4_2(4);
partial_p3_2(4) <= partial_p4_3(4);
HA_40 : HA port map(A=>partial_p4_0(5), B=>partial_p4_1(5), S=>partial_p3_1(5), C=>partial_p3_0(6));
partial_p3_2(5) <= partial_p4_2(5);
FA_364 : FA port map(A=>partial_p4_0(6), B=>partial_p4_1(6), Cin => partial_p4_2(6), S=>partial_p3_1(6), Cout=>partial_p3_0(7));
partial_p3_2(6) <= partial_p4_3(6);
FA_365 : FA port map(A=>partial_p4_0(7), B=>partial_p4_1(7), Cin => partial_p4_2(7), S=>partial_p3_1(7), Cout=>partial_p3_0(8));
partial_p3_2(7) <= partial_p4_3(7);
FA_366 : FA port map(A=>partial_p4_0(8), B=>partial_p4_1(8), Cin => partial_p4_2(8), S=>partial_p3_1(8), Cout=>partial_p3_0(9));
partial_p3_2(8) <= partial_p4_3(8);
FA_367 : FA port map(A=>partial_p4_0(9), B=>partial_p4_1(9), Cin => partial_p4_2(9), S=>partial_p3_1(9), Cout=>partial_p3_0(10));
partial_p3_2(9) <= partial_p4_3(9);
FA_368 : FA port map(A=>partial_p4_0(10), B=>partial_p4_1(10), Cin => partial_p4_2(10), S=>partial_p3_1(10), Cout=>partial_p3_0(11));
partial_p3_2(10) <= partial_p4_3(10);
FA_369 : FA port map(A=>partial_p4_0(11), B=>partial_p4_1(11), Cin => partial_p4_2(11), S=>partial_p3_1(11), Cout=>partial_p3_0(12));
partial_p3_2(11) <= partial_p4_3(11);
FA_370 : FA port map(A=>partial_p4_0(12), B=>partial_p4_1(12), Cin => partial_p4_2(12), S=>partial_p3_1(12), Cout=>partial_p3_0(13));
partial_p3_2(12) <= partial_p4_3(12);
FA_371 : FA port map(A=>partial_p4_0(13), B=>partial_p4_1(13), Cin => partial_p4_2(13), S=>partial_p3_1(13), Cout=>partial_p3_0(14));
partial_p3_2(13) <= partial_p4_3(13);
FA_372 : FA port map(A=>partial_p4_0(14), B=>partial_p4_1(14), Cin => partial_p4_2(14), S=>partial_p3_1(14), Cout=>partial_p3_0(15));
partial_p3_2(14) <= partial_p4_3(14);
FA_373 : FA port map(A=>partial_p4_0(15), B=>partial_p4_1(15), Cin => partial_p4_2(15), S=>partial_p3_1(15), Cout=>partial_p3_0(16));
partial_p3_2(15) <= partial_p4_3(15);
FA_374 : FA port map(A=>partial_p4_0(16), B=>partial_p4_1(16), Cin => partial_p4_2(16), S=>partial_p3_1(16), Cout=>partial_p3_0(17));
partial_p3_2(16) <= partial_p4_3(16);
FA_375 : FA port map(A=>partial_p4_0(17), B=>partial_p4_1(17), Cin => partial_p4_2(17), S=>partial_p3_1(17), Cout=>partial_p3_0(18));
partial_p3_2(17) <= partial_p4_3(17);
FA_376 : FA port map(A=>partial_p4_0(18), B=>partial_p4_1(18), Cin => partial_p4_2(18), S=>partial_p3_1(18), Cout=>partial_p3_0(19));
partial_p3_2(18) <= partial_p4_3(18);
FA_377 : FA port map(A=>partial_p4_0(19), B=>partial_p4_1(19), Cin => partial_p4_2(19), S=>partial_p3_1(19), Cout=>partial_p3_0(20));
partial_p3_2(19) <= partial_p4_3(19);
FA_378 : FA port map(A=>partial_p4_0(20), B=>partial_p4_1(20), Cin => partial_p4_2(20), S=>partial_p3_1(20), Cout=>partial_p3_0(21));
partial_p3_2(20) <= partial_p4_3(20);
FA_379 : FA port map(A=>partial_p4_0(21), B=>partial_p4_1(21), Cin => partial_p4_2(21), S=>partial_p3_1(21), Cout=>partial_p3_0(22));
partial_p3_2(21) <= partial_p4_3(21);
FA_380 : FA port map(A=>partial_p4_0(22), B=>partial_p4_1(22), Cin => partial_p4_2(22), S=>partial_p3_1(22), Cout=>partial_p3_0(23));
partial_p3_2(22) <= partial_p4_3(22);
FA_381 : FA port map(A=>partial_p4_0(23), B=>partial_p4_1(23), Cin => partial_p4_2(23), S=>partial_p3_1(23), Cout=>partial_p3_0(24));
partial_p3_2(23) <= partial_p4_3(23);
FA_382 : FA port map(A=>partial_p4_0(24), B=>partial_p4_1(24), Cin => partial_p4_2(24), S=>partial_p3_1(24), Cout=>partial_p3_0(25));
partial_p3_2(24) <= partial_p4_3(24);
FA_383 : FA port map(A=>partial_p4_0(25), B=>partial_p4_1(25), Cin => partial_p4_2(25), S=>partial_p3_1(25), Cout=>partial_p3_0(26));
partial_p3_2(25) <= partial_p4_3(25);
FA_384 : FA port map(A=>partial_p4_0(26), B=>partial_p4_1(26), Cin => partial_p4_2(26), S=>partial_p3_1(26), Cout=>partial_p3_0(27));
partial_p3_2(26) <= partial_p4_3(26);
FA_385 : FA port map(A=>partial_p4_0(27), B=>partial_p4_1(27), Cin => partial_p4_2(27), S=>partial_p3_1(27), Cout=>partial_p3_0(28));
partial_p3_2(27) <= partial_p4_3(27);
FA_386 : FA port map(A=>partial_p4_0(28), B=>partial_p4_1(28), Cin => partial_p4_2(28), S=>partial_p3_1(28), Cout=>partial_p3_0(29));
partial_p3_2(28) <= partial_p4_3(28);
FA_387 : FA port map(A=>partial_p4_0(29), B=>partial_p4_1(29), Cin => partial_p4_2(29), S=>partial_p3_1(29), Cout=>partial_p3_0(30));
partial_p3_2(29) <= partial_p4_3(29);
FA_388 : FA port map(A=>partial_p4_0(30), B=>partial_p4_1(30), Cin => partial_p4_2(30), S=>partial_p3_1(30), Cout=>partial_p3_0(31));
partial_p3_2(30) <= partial_p4_3(30);
FA_389 : FA port map(A=>partial_p4_0(31), B=>partial_p4_1(31), Cin => partial_p4_2(31), S=>partial_p3_1(31), Cout=>partial_p3_0(32));
partial_p3_2(31) <= partial_p4_3(31);
FA_390 : FA port map(A=>partial_p4_0(32), B=>partial_p4_1(32), Cin => partial_p4_2(32), S=>partial_p3_1(32), Cout=>partial_p3_0(33));
partial_p3_2(32) <= partial_p4_3(32);
FA_391 : FA port map(A=>partial_p4_0(33), B=>partial_p4_1(33), Cin => partial_p4_2(33), S=>partial_p3_1(33), Cout=>partial_p3_0(34));
partial_p3_2(33) <= partial_p4_3(33);
FA_392 : FA port map(A=>partial_p4_0(34), B=>partial_p4_1(34), Cin => partial_p4_2(34), S=>partial_p3_1(34), Cout=>partial_p3_0(35));
partial_p3_2(34) <= partial_p4_3(34);
FA_393 : FA port map(A=>partial_p4_0(35), B=>partial_p4_1(35), Cin => partial_p4_2(35), S=>partial_p3_1(35), Cout=>partial_p3_0(36));
partial_p3_2(35) <= partial_p4_3(35);
FA_394 : FA port map(A=>partial_p4_0(36), B=>partial_p4_1(36), Cin => partial_p4_2(36), S=>partial_p3_1(36), Cout=>partial_p3_0(37));
partial_p3_2(36) <= partial_p4_3(36);
FA_395 : FA port map(A=>partial_p4_0(37), B=>partial_p4_1(37), Cin => partial_p4_2(37), S=>partial_p3_1(37), Cout=>partial_p3_0(38));
partial_p3_2(37) <= partial_p4_3(37);
FA_396 : FA port map(A=>partial_p4_0(38), B=>partial_p4_1(38), Cin => partial_p4_2(38), S=>partial_p3_1(38), Cout=>partial_p3_0(39));
partial_p3_2(38) <= partial_p4_3(38);
FA_397 : FA port map(A=>partial_p4_0(39), B=>partial_p4_1(39), Cin => partial_p4_2(39), S=>partial_p3_1(39), Cout=>partial_p3_0(40));
partial_p3_2(39) <= partial_p4_3(39);
FA_398 : FA port map(A=>partial_p4_0(40), B=>partial_p4_1(40), Cin => partial_p4_2(40), S=>partial_p3_1(40), Cout=>partial_p3_0(41));
partial_p3_2(40) <= partial_p4_3(40);
FA_399 : FA port map(A=>partial_p4_0(41), B=>partial_p4_1(41), Cin => partial_p4_2(41), S=>partial_p3_1(41), Cout=>partial_p3_0(42));
partial_p3_2(41) <= partial_p4_3(41);
FA_400 : FA port map(A=>partial_p4_0(42), B=>partial_p4_1(42), Cin => partial_p4_2(42), S=>partial_p3_1(42), Cout=>partial_p3_0(43));
partial_p3_2(42) <= partial_p4_3(42);
FA_401 : FA port map(A=>partial_p4_0(43), B=>partial_p4_1(43), Cin => partial_p4_2(43), S=>partial_p3_1(43), Cout=>partial_p3_0(44));
partial_p3_2(43) <= partial_p4_3(43);
FA_402 : FA port map(A=>partial_p4_0(44), B=>partial_p4_1(44), Cin => partial_p4_2(44), S=>partial_p3_1(44), Cout=>partial_p3_0(45));
partial_p3_2(44) <= partial_p4_3(44);
FA_403 : FA port map(A=>partial_p4_0(45), B=>partial_p4_1(45), Cin => partial_p4_2(45), S=>partial_p3_1(45), Cout=>partial_p3_0(46));
partial_p3_2(45) <= partial_p4_3(45);
FA_404 : FA port map(A=>partial_p4_0(46), B=>partial_p4_1(46), Cin => partial_p4_2(46), S=>partial_p3_1(46), Cout=>partial_p3_0(47));
partial_p3_2(46) <= partial_p4_3(46);
FA_405 : FA port map(A=>partial_p4_0(47), B=>partial_p4_1(47), Cin => partial_p4_2(47), S=>partial_p3_1(47), Cout=>partial_p3_0(48));
partial_p3_2(47) <= partial_p4_3(47);
FA_406 : FA port map(A=>partial_p4_0(48), B=>partial_p4_1(48), Cin => partial_p4_2(48), S=>partial_p3_1(48), Cout=>partial_p3_0(49));
partial_p3_2(48) <= partial_p4_3(48);
FA_407 : FA port map(A=>partial_p4_0(49), B=>partial_p4_1(49), Cin => partial_p4_2(49), S=>partial_p3_1(49), Cout=>partial_p3_0(50));
partial_p3_2(49) <= partial_p4_3(49);
FA_408 : FA port map(A=>partial_p4_0(50), B=>partial_p4_1(50), Cin => partial_p4_2(50), S=>partial_p3_1(50), Cout=>partial_p3_0(51));
partial_p3_2(50) <= partial_p4_3(50);
FA_409 : FA port map(A=>partial_p4_0(51), B=>partial_p4_1(51), Cin => partial_p4_2(51), S=>partial_p3_1(51), Cout=>partial_p3_0(52));
partial_p3_2(51) <= partial_p4_3(51);
FA_410 : FA port map(A=>partial_p4_0(52), B=>partial_p4_1(52), Cin => partial_p4_2(52), S=>partial_p3_1(52), Cout=>partial_p3_0(53));
partial_p3_2(52) <= partial_p4_3(52);
FA_411 : FA port map(A=>partial_p4_0(53), B=>partial_p4_1(53), Cin => partial_p4_2(53), S=>partial_p3_1(53), Cout=>partial_p3_0(54));
partial_p3_2(53) <= partial_p4_3(53);
FA_412 : FA port map(A=>partial_p4_0(54), B=>partial_p4_1(54), Cin => partial_p4_2(54), S=>partial_p3_1(54), Cout=>partial_p3_0(55));
partial_p3_2(54) <= partial_p4_3(54);
FA_413 : FA port map(A=>partial_p4_0(55), B=>partial_p4_1(55), Cin => partial_p4_2(55), S=>partial_p3_1(55), Cout=>partial_p3_0(56));
partial_p3_2(55) <= partial_p4_3(55);
FA_414 : FA port map(A=>partial_p4_0(56), B=>partial_p4_1(56), Cin => partial_p4_2(56), S=>partial_p3_1(56), Cout=>partial_p3_0(57));
partial_p3_2(56) <= partial_p4_3(56);
FA_415 : FA port map(A=>partial_p4_0(57), B=>partial_p4_1(57), Cin => partial_p4_2(57), S=>partial_p3_1(57), Cout=>partial_p3_0(58));
partial_p3_2(57) <= partial_p4_3(57);
FA_416 : FA port map(A=>partial_p4_0(58), B=>partial_p4_1(58), Cin => partial_p4_2(58), S=>partial_p3_1(58), Cout=>partial_p3_0(59));
partial_p3_2(58) <= partial_p4_3(58);
FA_417 : FA port map(A=>partial_p4_0(59), B=>partial_p4_1(59), Cin => partial_p4_2(59), S=>partial_p3_1(59), Cout=>partial_p3_0(60));
partial_p3_2(59) <= partial_p4_3(59);
FA_418 : FA port map(A=>partial_p4_0(60), B=>partial_p4_1(60), Cin => partial_p4_2(60), S=>partial_p3_1(60), Cout=>partial_p3_0(61));
partial_p3_2(60) <= partial_p4_3(60);
FA_419 : FA port map(A=>partial_p4_0(61), B=>partial_p4_1(61), Cin => partial_p4_2(61), S=>partial_p3_1(61), Cout=>partial_p3_0(62));
partial_p3_2(61) <= partial_p4_3(61);
HA_41 : HA port map(A=>partial_p4_0(62), B=>partial_p4_1(62), S=>partial_p3_1(62), C=>partial_p3_0(63));
partial_p3_2(62) <= partial_p4_2(62);
partial_p3_1(63) <= partial_p4_0(63);
partial_p3_2(63) <= partial_p4_1(63);

--LEVEL 6

partial_p2_0(0) <= partial_p3_0(0);
partial_p2_1(0) <= partial_p3_1(0);
partial_p2_0(1) <= partial_p3_0(1);
partial_p2_1(1) <= partial_p3_1(1);
HA_42 : HA port map(A=>partial_p3_0(2), B=>partial_p3_1(2), S=>partial_p2_0(2), C=>partial_p2_0(3));
partial_p2_1(2) <= partial_p3_2(2);
HA_43 : HA port map(A=>partial_p3_0(3), B=>partial_p3_1(3), S=>partial_p2_1(3), C=>partial_p2_0(4));
FA_420 : FA port map(A=>partial_p3_0(4), B=>partial_p3_1(4), Cin => partial_p3_2(4), S=>partial_p2_1(4), Cout=>partial_p2_0(5));
FA_421 : FA port map(A=>partial_p3_0(5), B=>partial_p3_1(5), Cin => partial_p3_2(5), S=>partial_p2_1(5), Cout=>partial_p2_0(6));
FA_422 : FA port map(A=>partial_p3_0(6), B=>partial_p3_1(6), Cin => partial_p3_2(6), S=>partial_p2_1(6), Cout=>partial_p2_0(7));
FA_423 : FA port map(A=>partial_p3_0(7), B=>partial_p3_1(7), Cin => partial_p3_2(7), S=>partial_p2_1(7), Cout=>partial_p2_0(8));
FA_424 : FA port map(A=>partial_p3_0(8), B=>partial_p3_1(8), Cin => partial_p3_2(8), S=>partial_p2_1(8), Cout=>partial_p2_0(9));
FA_425 : FA port map(A=>partial_p3_0(9), B=>partial_p3_1(9), Cin => partial_p3_2(9), S=>partial_p2_1(9), Cout=>partial_p2_0(10));
FA_426 : FA port map(A=>partial_p3_0(10), B=>partial_p3_1(10), Cin => partial_p3_2(10), S=>partial_p2_1(10), Cout=>partial_p2_0(11));
FA_427 : FA port map(A=>partial_p3_0(11), B=>partial_p3_1(11), Cin => partial_p3_2(11), S=>partial_p2_1(11), Cout=>partial_p2_0(12));
FA_428 : FA port map(A=>partial_p3_0(12), B=>partial_p3_1(12), Cin => partial_p3_2(12), S=>partial_p2_1(12), Cout=>partial_p2_0(13));
FA_429 : FA port map(A=>partial_p3_0(13), B=>partial_p3_1(13), Cin => partial_p3_2(13), S=>partial_p2_1(13), Cout=>partial_p2_0(14));
FA_430 : FA port map(A=>partial_p3_0(14), B=>partial_p3_1(14), Cin => partial_p3_2(14), S=>partial_p2_1(14), Cout=>partial_p2_0(15));
FA_431 : FA port map(A=>partial_p3_0(15), B=>partial_p3_1(15), Cin => partial_p3_2(15), S=>partial_p2_1(15), Cout=>partial_p2_0(16));
FA_432 : FA port map(A=>partial_p3_0(16), B=>partial_p3_1(16), Cin => partial_p3_2(16), S=>partial_p2_1(16), Cout=>partial_p2_0(17));
FA_433 : FA port map(A=>partial_p3_0(17), B=>partial_p3_1(17), Cin => partial_p3_2(17), S=>partial_p2_1(17), Cout=>partial_p2_0(18));
FA_434 : FA port map(A=>partial_p3_0(18), B=>partial_p3_1(18), Cin => partial_p3_2(18), S=>partial_p2_1(18), Cout=>partial_p2_0(19));
FA_435 : FA port map(A=>partial_p3_0(19), B=>partial_p3_1(19), Cin => partial_p3_2(19), S=>partial_p2_1(19), Cout=>partial_p2_0(20));
FA_436 : FA port map(A=>partial_p3_0(20), B=>partial_p3_1(20), Cin => partial_p3_2(20), S=>partial_p2_1(20), Cout=>partial_p2_0(21));
FA_437 : FA port map(A=>partial_p3_0(21), B=>partial_p3_1(21), Cin => partial_p3_2(21), S=>partial_p2_1(21), Cout=>partial_p2_0(22));
FA_438 : FA port map(A=>partial_p3_0(22), B=>partial_p3_1(22), Cin => partial_p3_2(22), S=>partial_p2_1(22), Cout=>partial_p2_0(23));
FA_439 : FA port map(A=>partial_p3_0(23), B=>partial_p3_1(23), Cin => partial_p3_2(23), S=>partial_p2_1(23), Cout=>partial_p2_0(24));
FA_440 : FA port map(A=>partial_p3_0(24), B=>partial_p3_1(24), Cin => partial_p3_2(24), S=>partial_p2_1(24), Cout=>partial_p2_0(25));
FA_441 : FA port map(A=>partial_p3_0(25), B=>partial_p3_1(25), Cin => partial_p3_2(25), S=>partial_p2_1(25), Cout=>partial_p2_0(26));
FA_442 : FA port map(A=>partial_p3_0(26), B=>partial_p3_1(26), Cin => partial_p3_2(26), S=>partial_p2_1(26), Cout=>partial_p2_0(27));
FA_443 : FA port map(A=>partial_p3_0(27), B=>partial_p3_1(27), Cin => partial_p3_2(27), S=>partial_p2_1(27), Cout=>partial_p2_0(28));
FA_444 : FA port map(A=>partial_p3_0(28), B=>partial_p3_1(28), Cin => partial_p3_2(28), S=>partial_p2_1(28), Cout=>partial_p2_0(29));
FA_445 : FA port map(A=>partial_p3_0(29), B=>partial_p3_1(29), Cin => partial_p3_2(29), S=>partial_p2_1(29), Cout=>partial_p2_0(30));
FA_446 : FA port map(A=>partial_p3_0(30), B=>partial_p3_1(30), Cin => partial_p3_2(30), S=>partial_p2_1(30), Cout=>partial_p2_0(31));
FA_447 : FA port map(A=>partial_p3_0(31), B=>partial_p3_1(31), Cin => partial_p3_2(31), S=>partial_p2_1(31), Cout=>partial_p2_0(32));
FA_448 : FA port map(A=>partial_p3_0(32), B=>partial_p3_1(32), Cin => partial_p3_2(32), S=>partial_p2_1(32), Cout=>partial_p2_0(33));
FA_449 : FA port map(A=>partial_p3_0(33), B=>partial_p3_1(33), Cin => partial_p3_2(33), S=>partial_p2_1(33), Cout=>partial_p2_0(34));
FA_450 : FA port map(A=>partial_p3_0(34), B=>partial_p3_1(34), Cin => partial_p3_2(34), S=>partial_p2_1(34), Cout=>partial_p2_0(35));
FA_451 : FA port map(A=>partial_p3_0(35), B=>partial_p3_1(35), Cin => partial_p3_2(35), S=>partial_p2_1(35), Cout=>partial_p2_0(36));
FA_452 : FA port map(A=>partial_p3_0(36), B=>partial_p3_1(36), Cin => partial_p3_2(36), S=>partial_p2_1(36), Cout=>partial_p2_0(37));
FA_453 : FA port map(A=>partial_p3_0(37), B=>partial_p3_1(37), Cin => partial_p3_2(37), S=>partial_p2_1(37), Cout=>partial_p2_0(38));
FA_454 : FA port map(A=>partial_p3_0(38), B=>partial_p3_1(38), Cin => partial_p3_2(38), S=>partial_p2_1(38), Cout=>partial_p2_0(39));
FA_455 : FA port map(A=>partial_p3_0(39), B=>partial_p3_1(39), Cin => partial_p3_2(39), S=>partial_p2_1(39), Cout=>partial_p2_0(40));
FA_456 : FA port map(A=>partial_p3_0(40), B=>partial_p3_1(40), Cin => partial_p3_2(40), S=>partial_p2_1(40), Cout=>partial_p2_0(41));
FA_457 : FA port map(A=>partial_p3_0(41), B=>partial_p3_1(41), Cin => partial_p3_2(41), S=>partial_p2_1(41), Cout=>partial_p2_0(42));
FA_458 : FA port map(A=>partial_p3_0(42), B=>partial_p3_1(42), Cin => partial_p3_2(42), S=>partial_p2_1(42), Cout=>partial_p2_0(43));
FA_459 : FA port map(A=>partial_p3_0(43), B=>partial_p3_1(43), Cin => partial_p3_2(43), S=>partial_p2_1(43), Cout=>partial_p2_0(44));
FA_460 : FA port map(A=>partial_p3_0(44), B=>partial_p3_1(44), Cin => partial_p3_2(44), S=>partial_p2_1(44), Cout=>partial_p2_0(45));
FA_461 : FA port map(A=>partial_p3_0(45), B=>partial_p3_1(45), Cin => partial_p3_2(45), S=>partial_p2_1(45), Cout=>partial_p2_0(46));
FA_462 : FA port map(A=>partial_p3_0(46), B=>partial_p3_1(46), Cin => partial_p3_2(46), S=>partial_p2_1(46), Cout=>partial_p2_0(47));
FA_463 : FA port map(A=>partial_p3_0(47), B=>partial_p3_1(47), Cin => partial_p3_2(47), S=>partial_p2_1(47), Cout=>partial_p2_0(48));
FA_464 : FA port map(A=>partial_p3_0(48), B=>partial_p3_1(48), Cin => partial_p3_2(48), S=>partial_p2_1(48), Cout=>partial_p2_0(49));
FA_465 : FA port map(A=>partial_p3_0(49), B=>partial_p3_1(49), Cin => partial_p3_2(49), S=>partial_p2_1(49), Cout=>partial_p2_0(50));
FA_466 : FA port map(A=>partial_p3_0(50), B=>partial_p3_1(50), Cin => partial_p3_2(50), S=>partial_p2_1(50), Cout=>partial_p2_0(51));
FA_467 : FA port map(A=>partial_p3_0(51), B=>partial_p3_1(51), Cin => partial_p3_2(51), S=>partial_p2_1(51), Cout=>partial_p2_0(52));
FA_468 : FA port map(A=>partial_p3_0(52), B=>partial_p3_1(52), Cin => partial_p3_2(52), S=>partial_p2_1(52), Cout=>partial_p2_0(53));
FA_469 : FA port map(A=>partial_p3_0(53), B=>partial_p3_1(53), Cin => partial_p3_2(53), S=>partial_p2_1(53), Cout=>partial_p2_0(54));
FA_470 : FA port map(A=>partial_p3_0(54), B=>partial_p3_1(54), Cin => partial_p3_2(54), S=>partial_p2_1(54), Cout=>partial_p2_0(55));
FA_471 : FA port map(A=>partial_p3_0(55), B=>partial_p3_1(55), Cin => partial_p3_2(55), S=>partial_p2_1(55), Cout=>partial_p2_0(56));
FA_472 : FA port map(A=>partial_p3_0(56), B=>partial_p3_1(56), Cin => partial_p3_2(56), S=>partial_p2_1(56), Cout=>partial_p2_0(57));
FA_473 : FA port map(A=>partial_p3_0(57), B=>partial_p3_1(57), Cin => partial_p3_2(57), S=>partial_p2_1(57), Cout=>partial_p2_0(58));
FA_474 : FA port map(A=>partial_p3_0(58), B=>partial_p3_1(58), Cin => partial_p3_2(58), S=>partial_p2_1(58), Cout=>partial_p2_0(59));
FA_475 : FA port map(A=>partial_p3_0(59), B=>partial_p3_1(59), Cin => partial_p3_2(59), S=>partial_p2_1(59), Cout=>partial_p2_0(60));
FA_476 : FA port map(A=>partial_p3_0(60), B=>partial_p3_1(60), Cin => partial_p3_2(60), S=>partial_p2_1(60), Cout=>partial_p2_0(61));
FA_477 : FA port map(A=>partial_p3_0(61), B=>partial_p3_1(61), Cin => partial_p3_2(61), S=>partial_p2_1(61), Cout=>partial_p2_0(62));
FA_478 : FA port map(A=>partial_p3_0(62), B=>partial_p3_1(62), Cin => partial_p3_2(62), S=>partial_p2_1(62), Cout=>partial_p2_0(63));
FA_479 : FA port map(A=>partial_p3_0(63), B=>partial_p3_1(63), Cin => partial_p3_2(63), S=>partial_p2_1(63), Cout=>extra_carry);

product <= unsigned(partial_p2_0) + unsigned(partial_p2_1);

P <= std_logic_vector(product);

end beh;